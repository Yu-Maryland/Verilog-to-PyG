// Benchmark "Multi8" written by ABC on Sun Apr 16 09:24:28 2023

module Multi8 ( clock, 
    a0, a1, a2, a3, a4, a5, a6, a7, b0, b1, b2, b3, b4, b5, b6, b7,
    m00, m01, m02, m03, m04, m05, m06, m07, m08, m09, m10, m11, m12, m13,
    m14, m15  );
  input  clock;
  input  a0, a1, a2, a3, a4, a5, a6, a7, b0, b1, b2, b3, b4, b5, b6, b7;
  output m00, m01, m02, m03, m04, m05, m06, m07, m08, m09, m10, m11, m12, m13,
    m14, m15;
  reg n470_lo, n545_lo, n548_lo, n560_lo, n563_lo, n575_lo, n590_lo,
    n623_lo, n638_lo, n641_lo, n653_lo, n656_lo, n668_lo, n671_lo, n674_lo,
    n683_lo, n686_lo, n689_lo, n692_lo, n695_lo, n1001_o2, n996_o2,
    n1011_o2, n1056_o2, n1059_o2, n1074_o2, n1134_o2, n1135_o2, n1158_o2,
    n1237_o2, n1244_o2, n1266_o2, n1393_o2, n1394_o2, n1210_o2, n1211_o2,
    n1212_o2, n1437_o2, n1221_o2, n1230_o2, n1228_o2, n1229_o2, n1259_o2,
    n1265_o2, n1302_o2, n1326_o2, n1324_o2, n1325_o2, n1357_o2, n1648_o2,
    n1368_o2, n1654_o2, n1700_o2, n1448_o2, n1449_o2, n1490_o2, n1459_o2,
    n1460_o2, n1461_o2, n1464_o2, n1495_o2, n1496_o2, n1497_o2, n1605_o2,
    n1609_o2, n1520_o2, n1531_o2, n1670_o2, n467_o2, n466_o2, n1573_o2,
    n1606_o2, n1610_o2, n1625_o2, n662_lo_buf_o2, n468_o2, n519_o2,
    n1635_o2, n1682_o2, n371_o2, n370_o2, n520_o2, n1738_o2, n372_o2,
    n307_o2, n306_o2, n1719_o2, n1720_o2, n1721_o2, n1722_o2, n1743_o2,
    n523_o2, n567_o2, n308_o2, n1751_o2, n1752_o2, n1758_o2, n1765_o2,
    n527_lo_buf_o2, n677_lo_buf_o2, n606_o2, n657_o2, n568_o2,
    n647_lo_buf_o2, n542_lo_buf_o2, n617_lo_buf_o2, n335_o2, n287_o2,
    n530_o2, n334_o2, n286_o2, n557_lo_buf_o2, n288_o2, n638_1_o2, n673_o2,
    n415_o2, n672_o2, n571_o2, n646_o2, n414_o2, n608_o2, n659_o2, n637_o2,
    n461_o2, n551_o2, n618_o2, n336_o2, n367_o2, n572_lo_buf_o2, n304_o2,
    n509_o2, n591_o2, n525_o2, n615_o2, n416_o2, n402_o2, n489_o2, n533_o2,
    n463_o2, n553_o2, n620_o2, n508_o2, n590_1_o2, n368_o2, n482_lo_buf_o2,
    n497_lo_buf_o2, n587_lo_buf_o2, n602_lo_buf_o2, n659_lo_buf_o2,
    n446_o2, n536_o2, n375_o2, n474_o2, n426_o2, n351_o2, n632_lo_buf_o2,
    n404_o2, n491_o2, n445_o2, n535_o2, n467_lo_buf_o2, n328_o2, n387_o2,
    n305_o2, n340_o2, n423_o2, n274_o2, n275_o2, n428_o2, n353_o2, n327_o2,
    n386_o2, n512_lo_buf_o2, n281_o2, n533_lo_buf_o2, n608_lo_buf_o2,
    n293_o2, n292_o2, n276_o2, n524_lo_buf_o2, n283_o2;
  wire new_n577_, new_n579_, new_n581_1_, new_n583_, new_n585_, new_n587_,
    new_n589_, new_n591_1_, new_n593_, new_n596_1_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_1_, new_n602_, new_n603_, new_n605_,
    new_n606_1_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_1_,
    new_n612_, new_n613_, new_n614_, new_n616_1_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_1_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_1_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_1_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_1_,
    new_n637_, new_n638_, new_n639_, new_n641_1_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_1_, new_n647_, new_n648_, new_n649_,
    new_n652_, new_n653_, new_n655_, new_n656_1_, new_n657_, new_n660_,
    new_n661_1_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_1_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_1_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_1_, new_n678_, new_n680_,
    new_n682_, new_n688_, new_n689_, new_n690_, new_n691_1_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_1_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_1_, new_n702_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_1_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_1_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_1_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_1_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_1_, new_n732_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_1_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_1_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_1_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_1_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_1_,
    new_n762_, new_n765_, new_n766_1_, new_n768_, new_n769_, new_n771_1_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_1_, new_n777_,
    new_n779_, new_n780_, new_n781_1_, new_n782_, new_n783_, new_n784_,
    new_n786_1_, new_n787_, new_n788_, new_n795_, new_n796_1_, new_n798_,
    new_n799_, new_n800_, new_n801_1_, new_n802_, new_n804_, new_n805_,
    new_n806_1_, new_n807_, new_n809_, new_n810_, new_n811_1_, new_n813_,
    new_n815_, new_n816_1_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_1_, new_n822_, new_n823_, new_n825_, new_n826_1_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_1_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_1_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_1_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_1_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_1_,
    new_n852_, new_n854_, new_n855_, new_n856_1_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_1_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_1_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_1_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_1_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_1_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_1_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_1_, new_n897_, new_n898_, new_n901_1_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_1_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_1_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_1_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_1_,
    new_n922_, new_n923_, new_n925_, new_n926_1_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_1_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_1_, new_n940_, new_n941_1_, new_n942_, new_n943_,
    new_n944_, new_n946_1_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n953_, new_n954_, new_n955_, new_n956_1_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_1_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_1_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1007_, new_n1008_,
    new_n1009_, new_n1011_, new_n1012_, new_n1013_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1020_, new_n1021_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1045_, new_n1049_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1070_, new_n1071_, new_n1072_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1089_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1113_, new_n1114_,
    new_n1116_, new_n1117_, new_n1119_, new_n1121_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1129_, new_n1131_, new_n1136_,
    n66, n71, n76, n81, n86, n91, n96, n101, n106, n111, n116, n121, n126,
    n131, n136, n141, n146, n151, n156, n161, n166, n171, n176, n181, n186,
    n191, n196, n201, n206, n211, n216, n221, n226, n231, n236, n241, n246,
    n251, n256, n261, n266, n271, n276, n281, n286, n291, n296, n301, n306,
    n311, n316, n321, n326, n331, n336, n341, n346, n351, n356, n361, n366,
    n371, n376, n381, n386, n391, n396, n401, n406, n411, n416, n421, n426,
    n431, n436, n441, n446, n451, n456, n461, n466, n471, n476, n481, n486,
    n491, n496, n501, n506, n511, n516, n521, n526, n531, n536, n541, n546,
    n551, n556, n561, n566, n571, n576, n581, n586, n591, n596, n601, n606,
    n611, n616, n621, n626, n631, n636, n641, n646, n651, n656, n661, n666,
    n671, n676, n681, n686, n691, n696, n701, n706, n711, n716, n721, n726,
    n731, n736, n741, n746, n751, n756, n761, n766, n771, n776, n781, n786,
    n791, n796, n801, n806, n811, n816, n821, n826, n831, n836, n841, n846,
    n851, n856, n861, n866, n871, n876, n881, n886, n891, n896, n901, n906,
    n911, n916, n921, n926, n931, n936, n941, n946, n951, n956, n961, n966;
  AND2x2_ASAP7_75t_L        g000(.A(n470_lo), .B(n590_lo), .Y(m00));
  NOR2xp33_ASAP7_75t_L      g001(.A(n1001_o2), .B(n996_o2), .Y(new_n577_));
  NOR2xp33_ASAP7_75t_L      g002(.A(n1011_o2), .B(new_n577_), .Y(m01));
  NOR2xp33_ASAP7_75t_L      g003(.A(n1056_o2), .B(n1059_o2), .Y(new_n579_));
  NOR2xp33_ASAP7_75t_L      g004(.A(n1074_o2), .B(new_n579_), .Y(m02));
  NOR2xp33_ASAP7_75t_L      g005(.A(n1134_o2), .B(n1135_o2), .Y(new_n581_1_));
  NOR2xp33_ASAP7_75t_L      g006(.A(n1158_o2), .B(new_n581_1_), .Y(m03));
  NOR2xp33_ASAP7_75t_L      g007(.A(n1237_o2), .B(n1244_o2), .Y(new_n583_));
  NOR2xp33_ASAP7_75t_L      g008(.A(n1266_o2), .B(new_n583_), .Y(m04));
  NOR2xp33_ASAP7_75t_L      g009(.A(n1393_o2), .B(n1394_o2), .Y(new_n585_));
  NOR2xp33_ASAP7_75t_L      g010(.A(n1437_o2), .B(new_n585_), .Y(m05));
  NOR2xp33_ASAP7_75t_L      g011(.A(n1648_o2), .B(n1654_o2), .Y(new_n587_));
  NOR2xp33_ASAP7_75t_L      g012(.A(n1700_o2), .B(new_n587_), .Y(m06));
  NOR2xp33_ASAP7_75t_L      g013(.A(n467_o2), .B(n466_o2), .Y(new_n589_));
  NOR2xp33_ASAP7_75t_L      g014(.A(n468_o2), .B(new_n589_), .Y(m07));
  NOR2xp33_ASAP7_75t_L      g015(.A(n468_o2), .B(n519_o2), .Y(new_n591_1_));
  NOR2xp33_ASAP7_75t_L      g016(.A(n520_o2), .B(new_n591_1_), .Y(m08));
  INVx1_ASAP7_75t_L         g017(.A(n567_o2), .Y(new_n593_));
  AOI21xp33_ASAP7_75t_L     g018(.A1(new_n593_), .A2(n523_o2), .B(n568_o2), .Y(m09));
  XNOR2x2_ASAP7_75t_L       g019(.A(n571_o2), .B(n608_o2), .Y(m10));
  INVx1_ASAP7_75t_L         g020(.A(n571_o2), .Y(new_n596_1_));
  AOI21xp33_ASAP7_75t_L     g021(.A1(new_n596_1_), .A2(n608_o2), .B(n606_o2), .Y(new_n597_));
  INVx1_ASAP7_75t_L         g022(.A(n638_1_o2), .Y(new_n598_));
  INVx1_ASAP7_75t_L         g023(.A(n637_o2), .Y(new_n599_));
  NOR2xp33_ASAP7_75t_L      g024(.A(new_n598_), .B(new_n599_), .Y(new_n600_));
  INVx1_ASAP7_75t_L         g025(.A(new_n600_), .Y(new_n601_1_));
  NAND2xp33_ASAP7_75t_L     g026(.A(new_n598_), .B(new_n599_), .Y(new_n602_));
  NAND2xp33_ASAP7_75t_L     g027(.A(new_n602_), .B(new_n601_1_), .Y(new_n603_));
  XOR2x2_ASAP7_75t_L        g028(.A(new_n597_), .B(new_n603_), .Y(m11));
  INVx1_ASAP7_75t_L         g029(.A(n646_o2), .Y(new_n605_));
  NAND2xp33_ASAP7_75t_L     g030(.A(n659_o2), .B(new_n605_), .Y(new_n606_1_));
  INVx1_ASAP7_75t_L         g031(.A(n659_o2), .Y(new_n607_));
  NAND2xp33_ASAP7_75t_L     g032(.A(n646_o2), .B(new_n607_), .Y(new_n608_));
  NAND2xp33_ASAP7_75t_L     g033(.A(new_n606_1_), .B(new_n608_), .Y(new_n609_));
  NAND2xp33_ASAP7_75t_L     g034(.A(n545_lo), .B(n695_lo), .Y(new_n610_));
  XNOR2x2_ASAP7_75t_L       g035(.A(new_n610_), .B(new_n609_), .Y(new_n611_1_));
  O2A1O1Ixp33_ASAP7_75t_L   g036(.A1(new_n597_), .A2(new_n603_), .B(new_n601_1_), .C(new_n611_1_), .Y(new_n612_));
  A2O1A1O1Ixp25_ASAP7_75t_L g037(.A1(new_n596_1_), .A2(n608_o2), .B(n606_o2), .C(new_n602_), .D(new_n600_), .Y(new_n613_));
  AND2x2_ASAP7_75t_L        g038(.A(new_n611_1_), .B(new_n613_), .Y(new_n614_));
  NOR2xp33_ASAP7_75t_L      g039(.A(new_n612_), .B(new_n614_), .Y(m12));
  MAJIxp5_ASAP7_75t_L       g040(.A(new_n613_), .B(new_n610_), .C(new_n609_), .Y(new_n616_1_));
  INVx1_ASAP7_75t_L         g041(.A(n657_o2), .Y(new_n617_));
  NAND2xp33_ASAP7_75t_L     g042(.A(new_n617_), .B(new_n606_1_), .Y(new_n618_));
  INVx1_ASAP7_75t_L         g043(.A(n673_o2), .Y(new_n619_));
  NOR2xp33_ASAP7_75t_L      g044(.A(n672_o2), .B(new_n619_), .Y(new_n620_));
  INVx1_ASAP7_75t_L         g045(.A(n672_o2), .Y(new_n621_1_));
  NOR2xp33_ASAP7_75t_L      g046(.A(n673_o2), .B(new_n621_1_), .Y(new_n622_));
  NOR2xp33_ASAP7_75t_L      g047(.A(new_n620_), .B(new_n622_), .Y(new_n623_));
  NAND2xp33_ASAP7_75t_L     g048(.A(new_n618_), .B(new_n623_), .Y(new_n624_));
  NAND2xp33_ASAP7_75t_L     g049(.A(n673_o2), .B(new_n621_1_), .Y(new_n625_));
  NAND2xp33_ASAP7_75t_L     g050(.A(n672_o2), .B(new_n619_), .Y(new_n626_1_));
  NAND2xp33_ASAP7_75t_L     g051(.A(new_n625_), .B(new_n626_1_), .Y(new_n627_));
  NAND3xp33_ASAP7_75t_L     g052(.A(new_n627_), .B(new_n617_), .C(new_n606_1_), .Y(new_n628_));
  NAND2xp33_ASAP7_75t_L     g053(.A(n560_lo), .B(n695_lo), .Y(new_n629_));
  INVx1_ASAP7_75t_L         g054(.A(new_n629_), .Y(new_n630_));
  NAND3xp33_ASAP7_75t_L     g055(.A(new_n628_), .B(new_n624_), .C(new_n630_), .Y(new_n631_1_));
  O2A1O1Ixp33_ASAP7_75t_L   g056(.A1(n646_o2), .A2(new_n607_), .B(new_n617_), .C(new_n627_), .Y(new_n632_));
  NOR2xp33_ASAP7_75t_L      g057(.A(new_n618_), .B(new_n623_), .Y(new_n633_));
  OAI21xp33_ASAP7_75t_L     g058(.A1(new_n633_), .A2(new_n632_), .B(new_n629_), .Y(new_n634_));
  NAND3xp33_ASAP7_75t_L     g059(.A(new_n634_), .B(new_n631_1_), .C(new_n616_1_), .Y(new_n635_));
  MAJx2_ASAP7_75t_L         g060(.A(new_n609_), .B(new_n610_), .C(new_n613_), .Y(new_n636_1_));
  NOR3xp33_ASAP7_75t_L      g061(.A(new_n632_), .B(new_n633_), .C(new_n629_), .Y(new_n637_));
  AOI21xp33_ASAP7_75t_L     g062(.A1(new_n628_), .A2(new_n624_), .B(new_n630_), .Y(new_n638_));
  OAI21xp33_ASAP7_75t_L     g063(.A1(new_n638_), .A2(new_n637_), .B(new_n636_1_), .Y(new_n639_));
  AND2x2_ASAP7_75t_L        g064(.A(new_n639_), .B(new_n635_), .Y(m13));
  INVx1_ASAP7_75t_L         g065(.A(n575_lo), .Y(new_n641_1_));
  INVx1_ASAP7_75t_L         g066(.A(n695_lo), .Y(new_n642_));
  NOR2xp33_ASAP7_75t_L      g067(.A(new_n641_1_), .B(new_n642_), .Y(new_n643_));
  A2O1A1Ixp33_ASAP7_75t_L   g068(.A1(new_n618_), .A2(new_n626_1_), .B(new_n620_), .C(new_n643_), .Y(new_n644_));
  A2O1A1O1Ixp25_ASAP7_75t_L g069(.A1(new_n605_), .A2(n659_o2), .B(n657_o2), .C(new_n626_1_), .D(new_n620_), .Y(new_n645_));
  OAI21xp33_ASAP7_75t_L     g070(.A1(new_n641_1_), .A2(new_n642_), .B(new_n645_), .Y(new_n646_1_));
  NAND2xp33_ASAP7_75t_L     g071(.A(new_n644_), .B(new_n646_1_), .Y(new_n647_));
  O2A1O1Ixp33_ASAP7_75t_L   g072(.A1(new_n638_), .A2(new_n636_1_), .B(new_n631_1_), .C(new_n647_), .Y(new_n648_));
  AOI221xp5_ASAP7_75t_L     g073(.A1(new_n644_), .A2(new_n646_1_), .B1(new_n616_1_), .B2(new_n634_), .C(new_n637_), .Y(new_n649_));
  NOR2xp33_ASAP7_75t_L      g074(.A(new_n648_), .B(new_n649_), .Y(m14));
  A2O1A1Ixp33_ASAP7_75t_L   g075(.A1(new_n635_), .A2(new_n631_1_), .B(new_n647_), .C(new_n644_), .Y(m15));
  INVx1_ASAP7_75t_L         g076(.A(n692_lo), .Y(new_n652_));
  INVx1_ASAP7_75t_L         g077(.A(n1221_o2), .Y(new_n653_));
  NOR2xp33_ASAP7_75t_L      g078(.A(new_n652_), .B(new_n653_), .Y(n406));
  NAND2xp33_ASAP7_75t_L     g079(.A(n416_o2), .B(n463_o2), .Y(new_n655_));
  INVx1_ASAP7_75t_L         g080(.A(new_n655_), .Y(new_n656_1_));
  NOR2xp33_ASAP7_75t_L      g081(.A(n416_o2), .B(n463_o2), .Y(new_n657_));
  NOR2xp33_ASAP7_75t_L      g082(.A(new_n657_), .B(new_n656_1_), .Y(n411));
  NOR4xp25_ASAP7_75t_L      g083(.A(new_n656_1_), .B(new_n652_), .C(new_n653_), .D(new_n657_), .Y(n441));
  NAND2xp33_ASAP7_75t_L     g084(.A(n509_o2), .B(n508_o2), .Y(new_n660_));
  INVx1_ASAP7_75t_L         g085(.A(new_n660_), .Y(new_n661_1_));
  NOR2xp33_ASAP7_75t_L      g086(.A(n509_o2), .B(n508_o2), .Y(new_n662_));
  NOR2xp33_ASAP7_75t_L      g087(.A(new_n662_), .B(new_n661_1_), .Y(new_n663_));
  A2O1A1Ixp33_ASAP7_75t_L   g088(.A1(n416_o2), .A2(n463_o2), .B(n461_o2), .C(new_n663_), .Y(new_n664_));
  AOI21xp33_ASAP7_75t_L     g089(.A1(n416_o2), .A2(n463_o2), .B(n461_o2), .Y(new_n665_));
  INVx1_ASAP7_75t_L         g090(.A(new_n662_), .Y(new_n666_1_));
  NAND2xp33_ASAP7_75t_L     g091(.A(new_n660_), .B(new_n666_1_), .Y(new_n667_));
  NAND2xp33_ASAP7_75t_L     g092(.A(new_n665_), .B(new_n667_), .Y(new_n668_));
  NAND2xp33_ASAP7_75t_L     g093(.A(new_n668_), .B(new_n664_), .Y(new_n669_));
  NAND2xp33_ASAP7_75t_L     g094(.A(n692_lo), .B(n1210_o2), .Y(new_n670_));
  NOR2xp33_ASAP7_75t_L      g095(.A(new_n670_), .B(new_n669_), .Y(new_n671_1_));
  NOR2xp33_ASAP7_75t_L      g096(.A(new_n665_), .B(new_n667_), .Y(new_n672_));
  NOR3xp33_ASAP7_75t_L      g097(.A(new_n663_), .B(n461_o2), .C(new_n656_1_), .Y(new_n673_));
  NOR2xp33_ASAP7_75t_L      g098(.A(new_n672_), .B(new_n673_), .Y(new_n674_));
  INVx1_ASAP7_75t_L         g099(.A(new_n670_), .Y(new_n675_));
  NOR2xp33_ASAP7_75t_L      g100(.A(new_n675_), .B(new_n674_), .Y(new_n676_1_));
  NOR2xp33_ASAP7_75t_L      g101(.A(new_n671_1_), .B(new_n676_1_), .Y(n446));
  NAND2xp33_ASAP7_75t_L     g102(.A(n1464_o2), .B(n659_lo_buf_o2), .Y(new_n678_));
  INVx1_ASAP7_75t_L         g103(.A(new_n678_), .Y(n461));
  NOR2xp33_ASAP7_75t_L      g104(.A(n336_o2), .B(n367_o2), .Y(new_n680_));
  NOR2xp33_ASAP7_75t_L      g105(.A(n368_o2), .B(new_n680_), .Y(n466));
  INVx1_ASAP7_75t_L         g106(.A(n441), .Y(new_n682_));
  NOR3xp33_ASAP7_75t_L      g107(.A(new_n676_1_), .B(new_n671_1_), .C(new_n682_), .Y(n471));
  NOR3xp33_ASAP7_75t_L      g108(.A(new_n680_), .B(new_n678_), .C(n368_o2), .Y(n481));
  AND2x2_ASAP7_75t_L        g109(.A(n1743_o2), .B(n632_lo_buf_o2), .Y(n486));
  NOR2xp33_ASAP7_75t_L      g110(.A(n304_o2), .B(n305_o2), .Y(n491));
  MAJIxp5_ASAP7_75t_L       g111(.A(new_n674_), .B(n441), .C(new_n675_), .Y(n521));
  XOR2x2_ASAP7_75t_L        g112(.A(n525_o2), .B(n553_o2), .Y(new_n688_));
  NAND2xp33_ASAP7_75t_L     g113(.A(n1230_o2), .B(n677_lo_buf_o2), .Y(new_n689_));
  XNOR2x2_ASAP7_75t_L       g114(.A(new_n689_), .B(new_n688_), .Y(new_n690_));
  O2A1O1Ixp33_ASAP7_75t_L   g115(.A1(new_n665_), .A2(new_n667_), .B(new_n660_), .C(new_n690_), .Y(new_n691_1_));
  INVx1_ASAP7_75t_L         g116(.A(n461_o2), .Y(new_n692_));
  A2O1A1Ixp33_ASAP7_75t_L   g117(.A1(new_n655_), .A2(new_n692_), .B(new_n662_), .C(new_n660_), .Y(new_n693_));
  INVx1_ASAP7_75t_L         g118(.A(new_n689_), .Y(new_n694_));
  XNOR2x2_ASAP7_75t_L       g119(.A(new_n694_), .B(new_n688_), .Y(new_n695_));
  NOR2xp33_ASAP7_75t_L      g120(.A(new_n693_), .B(new_n695_), .Y(new_n696_1_));
  NAND2xp33_ASAP7_75t_L     g121(.A(n692_lo), .B(n1211_o2), .Y(new_n697_));
  NOR3xp33_ASAP7_75t_L      g122(.A(new_n691_1_), .B(new_n696_1_), .C(new_n697_), .Y(new_n698_));
  A2O1A1Ixp33_ASAP7_75t_L   g123(.A1(n509_o2), .A2(n508_o2), .B(new_n672_), .C(new_n695_), .Y(new_n699_));
  OA21x2_ASAP7_75t_L        g124(.A1(new_n662_), .A2(new_n665_), .B(new_n660_), .Y(new_n700_));
  NAND2xp33_ASAP7_75t_L     g125(.A(new_n700_), .B(new_n690_), .Y(new_n701_1_));
  AOI22xp33_ASAP7_75t_L     g126(.A1(n692_lo), .A2(n1211_o2), .B1(new_n701_1_), .B2(new_n699_), .Y(new_n702_));
  NOR2xp33_ASAP7_75t_L      g127(.A(new_n698_), .B(new_n702_), .Y(n526));
  NAND2xp33_ASAP7_75t_L     g128(.A(n1743_o2), .B(n632_lo_buf_o2), .Y(new_n704_));
  OR2x4_ASAP7_75t_L         g129(.A(n304_o2), .B(n305_o2), .Y(new_n705_));
  NOR2xp33_ASAP7_75t_L      g130(.A(new_n704_), .B(new_n705_), .Y(n531));
  NOR2xp33_ASAP7_75t_L      g131(.A(new_n689_), .B(new_n688_), .Y(new_n707_));
  NAND2xp33_ASAP7_75t_L     g132(.A(new_n689_), .B(new_n688_), .Y(new_n708_));
  AOI21xp33_ASAP7_75t_L     g133(.A1(new_n708_), .A2(new_n693_), .B(new_n707_), .Y(new_n709_));
  INVx1_ASAP7_75t_L         g134(.A(n525_o2), .Y(new_n710_));
  AOI21xp33_ASAP7_75t_L     g135(.A1(new_n710_), .A2(n553_o2), .B(n551_o2), .Y(new_n711_1_));
  XNOR2x2_ASAP7_75t_L       g136(.A(n591_o2), .B(n590_1_o2), .Y(new_n712_));
  NOR2xp33_ASAP7_75t_L      g137(.A(new_n711_1_), .B(new_n712_), .Y(new_n713_));
  INVx1_ASAP7_75t_L         g138(.A(n551_o2), .Y(new_n714_));
  INVx1_ASAP7_75t_L         g139(.A(n553_o2), .Y(new_n715_));
  OAI21xp33_ASAP7_75t_L     g140(.A1(n525_o2), .A2(new_n715_), .B(new_n714_), .Y(new_n716_1_));
  NAND2xp33_ASAP7_75t_L     g141(.A(n591_o2), .B(n590_1_o2), .Y(new_n717_));
  OR2x4_ASAP7_75t_L         g142(.A(n591_o2), .B(n590_1_o2), .Y(new_n718_));
  AOI21xp33_ASAP7_75t_L     g143(.A1(new_n717_), .A2(new_n718_), .B(new_n716_1_), .Y(new_n719_));
  INVx1_ASAP7_75t_L         g144(.A(n1265_o2), .Y(new_n720_));
  INVx1_ASAP7_75t_L         g145(.A(n677_lo_buf_o2), .Y(new_n721_1_));
  NOR2xp33_ASAP7_75t_L      g146(.A(new_n720_), .B(new_n721_1_), .Y(new_n722_));
  INVx1_ASAP7_75t_L         g147(.A(new_n722_), .Y(new_n723_));
  NOR3xp33_ASAP7_75t_L      g148(.A(new_n713_), .B(new_n719_), .C(new_n723_), .Y(new_n724_));
  NAND3xp33_ASAP7_75t_L     g149(.A(new_n716_1_), .B(new_n717_), .C(new_n718_), .Y(new_n725_));
  NAND2xp33_ASAP7_75t_L     g150(.A(new_n711_1_), .B(new_n712_), .Y(new_n726_1_));
  AOI21xp33_ASAP7_75t_L     g151(.A1(new_n725_), .A2(new_n726_1_), .B(new_n722_), .Y(new_n727_));
  NOR3xp33_ASAP7_75t_L      g152(.A(new_n724_), .B(new_n727_), .C(new_n709_), .Y(new_n728_));
  MAJIxp5_ASAP7_75t_L       g153(.A(new_n700_), .B(new_n689_), .C(new_n688_), .Y(new_n729_));
  NAND3xp33_ASAP7_75t_L     g154(.A(new_n725_), .B(new_n726_1_), .C(new_n722_), .Y(new_n730_));
  OAI21xp33_ASAP7_75t_L     g155(.A1(new_n719_), .A2(new_n713_), .B(new_n723_), .Y(new_n731_1_));
  AOI21xp33_ASAP7_75t_L     g156(.A1(new_n730_), .A2(new_n731_1_), .B(new_n729_), .Y(new_n732_));
  INVx1_ASAP7_75t_L         g157(.A(n1230_o2), .Y(new_n733_));
  NOR2xp33_ASAP7_75t_L      g158(.A(new_n652_), .B(new_n733_), .Y(new_n734_));
  INVx1_ASAP7_75t_L         g159(.A(new_n734_), .Y(new_n735_));
  NOR3xp33_ASAP7_75t_L      g160(.A(new_n728_), .B(new_n732_), .C(new_n735_), .Y(n566));
  INVx1_ASAP7_75t_L         g161(.A(n615_o2), .Y(new_n737_));
  NAND2xp33_ASAP7_75t_L     g162(.A(n620_o2), .B(new_n737_), .Y(new_n738_));
  INVx1_ASAP7_75t_L         g163(.A(n620_o2), .Y(new_n739_));
  NAND2xp33_ASAP7_75t_L     g164(.A(n615_o2), .B(new_n739_), .Y(new_n740_));
  AND2x2_ASAP7_75t_L        g165(.A(n1326_o2), .B(n662_lo_buf_o2), .Y(new_n741_1_));
  NAND3xp33_ASAP7_75t_L     g166(.A(new_n738_), .B(new_n740_), .C(new_n741_1_), .Y(new_n742_));
  INVx1_ASAP7_75t_L         g167(.A(new_n717_), .Y(new_n743_));
  A2O1A1O1Ixp25_ASAP7_75t_L g168(.A1(new_n710_), .A2(n553_o2), .B(n551_o2), .C(new_n718_), .D(new_n743_), .Y(new_n744_));
  AOI21xp33_ASAP7_75t_L     g169(.A1(new_n738_), .A2(new_n740_), .B(new_n741_1_), .Y(new_n745_));
  INVx1_ASAP7_75t_L         g170(.A(n618_o2), .Y(new_n746_1_));
  NAND2xp33_ASAP7_75t_L     g171(.A(n1368_o2), .B(n662_lo_buf_o2), .Y(new_n747_));
  O2A1O1Ixp33_ASAP7_75t_L   g172(.A1(n615_o2), .A2(new_n739_), .B(new_n746_1_), .C(new_n747_), .Y(new_n748_));
  AOI221xp5_ASAP7_75t_L     g173(.A1(n1368_o2), .A2(n662_lo_buf_o2), .B1(n620_o2), .B2(new_n737_), .C(n618_o2), .Y(new_n749_));
  OR2x4_ASAP7_75t_L         g174(.A(new_n748_), .B(new_n749_), .Y(new_n750_));
  O2A1O1Ixp33_ASAP7_75t_L   g175(.A1(new_n744_), .A2(new_n745_), .B(new_n742_), .C(new_n750_), .Y(new_n751_1_));
  NOR2xp33_ASAP7_75t_L      g176(.A(n615_o2), .B(new_n739_), .Y(new_n752_));
  NOR2xp33_ASAP7_75t_L      g177(.A(n620_o2), .B(new_n737_), .Y(new_n753_));
  NAND2xp33_ASAP7_75t_L     g178(.A(n1326_o2), .B(n662_lo_buf_o2), .Y(new_n754_));
  NOR3xp33_ASAP7_75t_L      g179(.A(new_n752_), .B(new_n753_), .C(new_n754_), .Y(new_n755_));
  NAND2xp33_ASAP7_75t_L     g180(.A(n553_o2), .B(new_n710_), .Y(new_n756_1_));
  NOR2xp33_ASAP7_75t_L      g181(.A(n591_o2), .B(n590_1_o2), .Y(new_n757_));
  A2O1A1Ixp33_ASAP7_75t_L   g182(.A1(new_n756_1_), .A2(new_n714_), .B(new_n757_), .C(new_n717_), .Y(new_n758_));
  OAI21xp33_ASAP7_75t_L     g183(.A1(new_n752_), .A2(new_n753_), .B(new_n754_), .Y(new_n759_));
  NOR2xp33_ASAP7_75t_L      g184(.A(new_n748_), .B(new_n749_), .Y(new_n760_));
  AOI211xp5_ASAP7_75t_L     g185(.A1(new_n758_), .A2(new_n759_), .B(new_n755_), .C(new_n760_), .Y(new_n761_1_));
  NAND2xp33_ASAP7_75t_L     g186(.A(n1326_o2), .B(n677_lo_buf_o2), .Y(new_n762_));
  NOR3xp33_ASAP7_75t_L      g187(.A(new_n751_1_), .B(new_n761_1_), .C(new_n762_), .Y(n571));
  NOR3xp33_ASAP7_75t_L      g188(.A(new_n702_), .B(new_n698_), .C(n521), .Y(n576));
  INVx1_ASAP7_75t_L         g189(.A(n641_lo), .Y(new_n765_));
  INVx1_ASAP7_75t_L         g190(.A(n1743_o2), .Y(new_n766_1_));
  NOR2xp33_ASAP7_75t_L      g191(.A(new_n765_), .B(new_n766_1_), .Y(n596));
  INVx1_ASAP7_75t_L         g192(.A(n467_lo_buf_o2), .Y(new_n768_));
  INVx1_ASAP7_75t_L         g193(.A(n608_lo_buf_o2), .Y(new_n769_));
  NOR2xp33_ASAP7_75t_L      g194(.A(new_n768_), .B(new_n769_), .Y(n601));
  INVx1_ASAP7_75t_L         g195(.A(n426_o2), .Y(new_n771_1_));
  INVx1_ASAP7_75t_L         g196(.A(n428_o2), .Y(new_n772_));
  NAND2xp33_ASAP7_75t_L     g197(.A(n1722_o2), .B(n572_lo_buf_o2), .Y(new_n773_));
  O2A1O1Ixp33_ASAP7_75t_L   g198(.A1(n423_o2), .A2(new_n772_), .B(new_n771_1_), .C(new_n773_), .Y(new_n774_));
  INVx1_ASAP7_75t_L         g199(.A(n617_lo_buf_o2), .Y(new_n775_));
  INVx1_ASAP7_75t_L         g200(.A(n572_lo_buf_o2), .Y(new_n776_1_));
  NOR2xp33_ASAP7_75t_L      g201(.A(new_n775_), .B(new_n776_1_), .Y(new_n777_));
  AND2x2_ASAP7_75t_L        g202(.A(new_n774_), .B(new_n777_), .Y(n606));
  AND2x2_ASAP7_75t_L        g203(.A(n328_o2), .B(n327_o2), .Y(new_n779_));
  NOR2xp33_ASAP7_75t_L      g204(.A(n328_o2), .B(n327_o2), .Y(new_n780_));
  NOR4xp25_ASAP7_75t_L      g205(.A(new_n705_), .B(new_n704_), .C(new_n779_), .D(new_n780_), .Y(new_n781_1_));
  NAND2xp33_ASAP7_75t_L     g206(.A(n328_o2), .B(n327_o2), .Y(new_n782_));
  OR2x4_ASAP7_75t_L         g207(.A(n328_o2), .B(n327_o2), .Y(new_n783_));
  AOI21xp33_ASAP7_75t_L     g208(.A1(new_n782_), .A2(new_n783_), .B(n531), .Y(new_n784_));
  NOR2xp33_ASAP7_75t_L      g209(.A(new_n781_1_), .B(new_n784_), .Y(n611));
  NAND2xp33_ASAP7_75t_L     g210(.A(n276_o2), .B(n283_o2), .Y(new_n786_1_));
  INVx1_ASAP7_75t_L         g211(.A(new_n786_1_), .Y(new_n787_));
  NOR2xp33_ASAP7_75t_L      g212(.A(n276_o2), .B(n283_o2), .Y(new_n788_));
  NOR2xp33_ASAP7_75t_L      g213(.A(new_n788_), .B(new_n787_), .Y(n616));
  NOR4xp25_ASAP7_75t_L      g214(.A(new_n787_), .B(new_n768_), .C(new_n769_), .D(new_n788_), .Y(n626));
  NOR2xp33_ASAP7_75t_L      g215(.A(new_n652_), .B(new_n720_), .Y(n631));
  AND2x2_ASAP7_75t_L        g216(.A(n1368_o2), .B(n677_lo_buf_o2), .Y(n636));
  AND2x2_ASAP7_75t_L        g217(.A(n674_lo), .B(n1464_o2), .Y(n641));
  A2O1A1O1Ixp25_ASAP7_75t_L g218(.A1(new_n759_), .A2(new_n758_), .B(new_n755_), .C(new_n760_), .D(new_n748_), .Y(n646));
  MAJIxp5_ASAP7_75t_L       g219(.A(new_n669_), .B(new_n682_), .C(new_n670_), .Y(new_n795_));
  OAI21xp33_ASAP7_75t_L     g220(.A1(new_n696_1_), .A2(new_n691_1_), .B(new_n697_), .Y(new_n796_1_));
  AOI21xp33_ASAP7_75t_L     g221(.A1(new_n796_1_), .A2(new_n795_), .B(new_n698_), .Y(n651));
  NOR3xp33_ASAP7_75t_L      g222(.A(new_n744_), .B(new_n755_), .C(new_n745_), .Y(new_n798_));
  AOI21xp33_ASAP7_75t_L     g223(.A1(new_n759_), .A2(new_n742_), .B(new_n758_), .Y(new_n799_));
  NAND2xp33_ASAP7_75t_L     g224(.A(n1302_o2), .B(n677_lo_buf_o2), .Y(new_n800_));
  NOR3xp33_ASAP7_75t_L      g225(.A(new_n798_), .B(new_n799_), .C(new_n800_), .Y(new_n801_1_));
  OAI21xp33_ASAP7_75t_L     g226(.A1(new_n799_), .A2(new_n798_), .B(new_n800_), .Y(new_n802_));
  A2O1A1O1Ixp25_ASAP7_75t_L g227(.A1(new_n729_), .A2(new_n731_1_), .B(new_n724_), .C(new_n802_), .D(new_n801_1_), .Y(n656));
  XNOR2x2_ASAP7_75t_L       g228(.A(n375_o2), .B(n404_o2), .Y(new_n804_));
  NAND2xp33_ASAP7_75t_L     g229(.A(n1459_o2), .B(n659_lo_buf_o2), .Y(new_n805_));
  INVx1_ASAP7_75t_L         g230(.A(new_n805_), .Y(new_n806_1_));
  XNOR2x2_ASAP7_75t_L       g231(.A(new_n806_1_), .B(new_n804_), .Y(new_n807_));
  XNOR2x2_ASAP7_75t_L       g232(.A(n481), .B(new_n807_), .Y(n661));
  NAND3xp33_ASAP7_75t_L     g233(.A(new_n730_), .B(new_n731_1_), .C(new_n729_), .Y(new_n809_));
  OAI21xp33_ASAP7_75t_L     g234(.A1(new_n727_), .A2(new_n724_), .B(new_n709_), .Y(new_n810_));
  AOI21xp33_ASAP7_75t_L     g235(.A1(new_n810_), .A2(new_n809_), .B(new_n734_), .Y(new_n811_1_));
  NOR2xp33_ASAP7_75t_L      g236(.A(new_n811_1_), .B(n566), .Y(n666));
  OA21x2_ASAP7_75t_L        g237(.A1(new_n761_1_), .A2(new_n751_1_), .B(new_n762_), .Y(new_n813_));
  NOR2xp33_ASAP7_75t_L      g238(.A(n571), .B(new_n813_), .Y(n671));
  AOI21xp33_ASAP7_75t_L     g239(.A1(new_n729_), .A2(new_n731_1_), .B(new_n724_), .Y(new_n815_));
  NAND3xp33_ASAP7_75t_L     g240(.A(new_n758_), .B(new_n759_), .C(new_n742_), .Y(new_n816_1_));
  OAI21xp33_ASAP7_75t_L     g241(.A1(new_n745_), .A2(new_n755_), .B(new_n744_), .Y(new_n817_));
  INVx1_ASAP7_75t_L         g242(.A(new_n800_), .Y(new_n818_));
  AOI21xp33_ASAP7_75t_L     g243(.A1(new_n816_1_), .A2(new_n817_), .B(new_n818_), .Y(new_n819_));
  NOR3xp33_ASAP7_75t_L      g244(.A(new_n801_1_), .B(new_n819_), .C(new_n815_), .Y(new_n820_));
  NAND3xp33_ASAP7_75t_L     g245(.A(new_n816_1_), .B(new_n817_), .C(new_n818_), .Y(new_n821_1_));
  OAI21xp33_ASAP7_75t_L     g246(.A1(new_n709_), .A2(new_n727_), .B(new_n730_), .Y(new_n822_));
  AOI21xp33_ASAP7_75t_L     g247(.A1(new_n802_), .A2(new_n821_1_), .B(new_n822_), .Y(new_n823_));
  NOR2xp33_ASAP7_75t_L      g248(.A(new_n823_), .B(new_n820_), .Y(n676));
  MAJIxp5_ASAP7_75t_L       g249(.A(n481), .B(new_n806_1_), .C(new_n804_), .Y(new_n825_));
  INVx1_ASAP7_75t_L         g250(.A(n375_o2), .Y(new_n826_1_));
  AOI21xp33_ASAP7_75t_L     g251(.A1(new_n826_1_), .A2(n404_o2), .B(n402_o2), .Y(new_n827_));
  XNOR2x2_ASAP7_75t_L       g252(.A(n446_o2), .B(n445_o2), .Y(new_n828_));
  NOR2xp33_ASAP7_75t_L      g253(.A(new_n827_), .B(new_n828_), .Y(new_n829_));
  INVx1_ASAP7_75t_L         g254(.A(n402_o2), .Y(new_n830_));
  INVx1_ASAP7_75t_L         g255(.A(n404_o2), .Y(new_n831_1_));
  OAI21xp33_ASAP7_75t_L     g256(.A1(n375_o2), .A2(new_n831_1_), .B(new_n830_), .Y(new_n832_));
  NAND2xp33_ASAP7_75t_L     g257(.A(n446_o2), .B(n445_o2), .Y(new_n833_));
  OR2x4_ASAP7_75t_L         g258(.A(n446_o2), .B(n445_o2), .Y(new_n834_));
  AOI21xp33_ASAP7_75t_L     g259(.A1(new_n833_), .A2(new_n834_), .B(new_n832_), .Y(new_n835_));
  INVx1_ASAP7_75t_L         g260(.A(n1460_o2), .Y(new_n836_1_));
  INVx1_ASAP7_75t_L         g261(.A(n659_lo_buf_o2), .Y(new_n837_));
  NOR2xp33_ASAP7_75t_L      g262(.A(new_n836_1_), .B(new_n837_), .Y(new_n838_));
  INVx1_ASAP7_75t_L         g263(.A(new_n838_), .Y(new_n839_));
  NOR3xp33_ASAP7_75t_L      g264(.A(new_n829_), .B(new_n835_), .C(new_n839_), .Y(new_n840_));
  NAND3xp33_ASAP7_75t_L     g265(.A(new_n832_), .B(new_n833_), .C(new_n834_), .Y(new_n841_1_));
  NAND2xp33_ASAP7_75t_L     g266(.A(new_n827_), .B(new_n828_), .Y(new_n842_));
  AOI21xp33_ASAP7_75t_L     g267(.A1(new_n841_1_), .A2(new_n842_), .B(new_n838_), .Y(new_n843_));
  NOR3xp33_ASAP7_75t_L      g268(.A(new_n840_), .B(new_n843_), .C(new_n825_), .Y(new_n844_));
  MAJx2_ASAP7_75t_L         g269(.A(new_n804_), .B(new_n806_1_), .C(n481), .Y(new_n845_));
  NAND3xp33_ASAP7_75t_L     g270(.A(new_n841_1_), .B(new_n842_), .C(new_n838_), .Y(new_n846_1_));
  OAI21xp33_ASAP7_75t_L     g271(.A1(new_n835_), .A2(new_n829_), .B(new_n839_), .Y(new_n847_));
  AOI21xp33_ASAP7_75t_L     g272(.A1(new_n846_1_), .A2(new_n847_), .B(new_n845_), .Y(new_n848_));
  INVx1_ASAP7_75t_L         g273(.A(n674_lo), .Y(new_n849_));
  INVx1_ASAP7_75t_L         g274(.A(n1459_o2), .Y(new_n850_));
  NOR2xp33_ASAP7_75t_L      g275(.A(new_n849_), .B(new_n850_), .Y(new_n851_1_));
  INVx1_ASAP7_75t_L         g276(.A(new_n851_1_), .Y(new_n852_));
  NOR3xp33_ASAP7_75t_L      g277(.A(new_n844_), .B(new_n848_), .C(new_n852_), .Y(n681));
  XOR2x2_ASAP7_75t_L        g278(.A(n474_o2), .B(n491_o2), .Y(new_n854_));
  NAND2xp33_ASAP7_75t_L     g279(.A(n1531_o2), .B(n647_lo_buf_o2), .Y(new_n855_));
  NOR2xp33_ASAP7_75t_L      g280(.A(new_n855_), .B(new_n854_), .Y(new_n856_1_));
  NOR2xp33_ASAP7_75t_L      g281(.A(n446_o2), .B(n445_o2), .Y(new_n857_));
  OAI21xp33_ASAP7_75t_L     g282(.A1(new_n857_), .A2(new_n827_), .B(new_n833_), .Y(new_n858_));
  NAND2xp33_ASAP7_75t_L     g283(.A(new_n855_), .B(new_n854_), .Y(new_n859_));
  AOI21xp33_ASAP7_75t_L     g284(.A1(new_n858_), .A2(new_n859_), .B(new_n856_1_), .Y(new_n860_));
  INVx1_ASAP7_75t_L         g285(.A(n474_o2), .Y(new_n861_1_));
  AOI21xp33_ASAP7_75t_L     g286(.A1(new_n861_1_), .A2(n491_o2), .B(n489_o2), .Y(new_n862_));
  AND2x2_ASAP7_75t_L        g287(.A(n536_o2), .B(n535_o2), .Y(new_n863_));
  NOR2xp33_ASAP7_75t_L      g288(.A(n536_o2), .B(n535_o2), .Y(new_n864_));
  NOR3xp33_ASAP7_75t_L      g289(.A(new_n862_), .B(new_n863_), .C(new_n864_), .Y(new_n865_));
  INVx1_ASAP7_75t_L         g290(.A(n489_o2), .Y(new_n866_1_));
  INVx1_ASAP7_75t_L         g291(.A(n491_o2), .Y(new_n867_));
  OAI21xp33_ASAP7_75t_L     g292(.A1(n474_o2), .A2(new_n867_), .B(new_n866_1_), .Y(new_n868_));
  NAND2xp33_ASAP7_75t_L     g293(.A(n536_o2), .B(n535_o2), .Y(new_n869_));
  OR2x4_ASAP7_75t_L         g294(.A(n536_o2), .B(n535_o2), .Y(new_n870_));
  AOI21xp33_ASAP7_75t_L     g295(.A1(new_n869_), .A2(new_n870_), .B(new_n868_), .Y(new_n871_1_));
  NAND2xp33_ASAP7_75t_L     g296(.A(n1573_o2), .B(n647_lo_buf_o2), .Y(new_n872_));
  NOR3xp33_ASAP7_75t_L      g297(.A(new_n865_), .B(new_n871_1_), .C(new_n872_), .Y(new_n873_));
  NAND3xp33_ASAP7_75t_L     g298(.A(new_n868_), .B(new_n870_), .C(new_n869_), .Y(new_n874_));
  OAI21xp33_ASAP7_75t_L     g299(.A1(new_n863_), .A2(new_n864_), .B(new_n862_), .Y(new_n875_));
  INVx1_ASAP7_75t_L         g300(.A(new_n872_), .Y(new_n876_1_));
  AOI21xp33_ASAP7_75t_L     g301(.A1(new_n874_), .A2(new_n875_), .B(new_n876_1_), .Y(new_n877_));
  NOR3xp33_ASAP7_75t_L      g302(.A(new_n873_), .B(new_n860_), .C(new_n877_), .Y(new_n878_));
  NAND2xp33_ASAP7_75t_L     g303(.A(n491_o2), .B(new_n861_1_), .Y(new_n879_));
  NAND2xp33_ASAP7_75t_L     g304(.A(n474_o2), .B(new_n867_), .Y(new_n880_));
  AND2x2_ASAP7_75t_L        g305(.A(n1531_o2), .B(n647_lo_buf_o2), .Y(new_n881_1_));
  NAND3xp33_ASAP7_75t_L     g306(.A(new_n879_), .B(new_n880_), .C(new_n881_1_), .Y(new_n882_));
  AND2x2_ASAP7_75t_L        g307(.A(n446_o2), .B(n445_o2), .Y(new_n883_));
  A2O1A1O1Ixp25_ASAP7_75t_L g308(.A1(new_n826_1_), .A2(n404_o2), .B(n402_o2), .C(new_n834_), .D(new_n883_), .Y(new_n884_));
  AOI21xp33_ASAP7_75t_L     g309(.A1(new_n879_), .A2(new_n880_), .B(new_n881_1_), .Y(new_n885_));
  OAI21xp33_ASAP7_75t_L     g310(.A1(new_n885_), .A2(new_n884_), .B(new_n882_), .Y(new_n886_1_));
  NAND3xp33_ASAP7_75t_L     g311(.A(new_n874_), .B(new_n875_), .C(new_n876_1_), .Y(new_n887_));
  OAI21xp33_ASAP7_75t_L     g312(.A1(new_n871_1_), .A2(new_n865_), .B(new_n872_), .Y(new_n888_));
  AOI21xp33_ASAP7_75t_L     g313(.A1(new_n888_), .A2(new_n887_), .B(new_n886_1_), .Y(new_n889_));
  NAND2xp33_ASAP7_75t_L     g314(.A(n1531_o2), .B(n659_lo_buf_o2), .Y(new_n890_));
  NOR3xp33_ASAP7_75t_L      g315(.A(new_n878_), .B(new_n889_), .C(new_n890_), .Y(n686));
  OAI211xp5_ASAP7_75t_L     g316(.A1(n530_o2), .A2(n533_o2), .B(n1682_o2), .C(n1738_o2), .Y(new_n892_));
  A2O1A1O1Ixp25_ASAP7_75t_L g317(.A1(new_n861_1_), .A2(n491_o2), .B(n489_o2), .C(new_n870_), .D(new_n863_), .Y(new_n893_));
  NOR2xp33_ASAP7_75t_L      g318(.A(n530_o2), .B(n533_o2), .Y(new_n894_));
  NAND2xp33_ASAP7_75t_L     g319(.A(n1682_o2), .B(n1738_o2), .Y(new_n895_));
  NAND2xp33_ASAP7_75t_L     g320(.A(new_n895_), .B(new_n894_), .Y(new_n896_1_));
  NAND2xp33_ASAP7_75t_L     g321(.A(new_n892_), .B(new_n896_1_), .Y(new_n897_));
  NAND2xp33_ASAP7_75t_L     g322(.A(n1682_o2), .B(n647_lo_buf_o2), .Y(new_n898_));
  O2A1O1Ixp33_ASAP7_75t_L   g323(.A1(new_n897_), .A2(new_n893_), .B(new_n892_), .C(new_n898_), .Y(n691));
  NOR4xp25_ASAP7_75t_L      g324(.A(new_n784_), .B(new_n765_), .C(new_n766_1_), .D(new_n781_1_), .Y(n696));
  INVx1_ASAP7_75t_L         g325(.A(n1719_o2), .Y(new_n901_1_));
  AOI31xp33_ASAP7_75t_L     g326(.A1(new_n783_), .A2(n486), .A3(n491), .B(new_n779_), .Y(new_n902_));
  INVx1_ASAP7_75t_L         g327(.A(n340_o2), .Y(new_n903_));
  NAND2xp33_ASAP7_75t_L     g328(.A(n353_o2), .B(new_n903_), .Y(new_n904_));
  INVx1_ASAP7_75t_L         g329(.A(n353_o2), .Y(new_n905_));
  NAND2xp33_ASAP7_75t_L     g330(.A(n340_o2), .B(new_n905_), .Y(new_n906_1_));
  NAND2xp33_ASAP7_75t_L     g331(.A(n1720_o2), .B(n632_lo_buf_o2), .Y(new_n907_));
  INVx1_ASAP7_75t_L         g332(.A(new_n907_), .Y(new_n908_));
  NAND3xp33_ASAP7_75t_L     g333(.A(new_n908_), .B(new_n904_), .C(new_n906_1_), .Y(new_n909_));
  XOR2x2_ASAP7_75t_L        g334(.A(n340_o2), .B(n353_o2), .Y(new_n910_));
  NAND2xp33_ASAP7_75t_L     g335(.A(new_n907_), .B(new_n910_), .Y(new_n911_1_));
  NAND2xp33_ASAP7_75t_L     g336(.A(new_n911_1_), .B(new_n909_), .Y(new_n912_));
  NOR2xp33_ASAP7_75t_L      g337(.A(new_n902_), .B(new_n912_), .Y(new_n913_));
  OAI31xp33_ASAP7_75t_L     g338(.A1(new_n705_), .A2(new_n704_), .A3(new_n780_), .B(new_n782_), .Y(new_n914_));
  NOR2xp33_ASAP7_75t_L      g339(.A(new_n907_), .B(new_n910_), .Y(new_n915_));
  AOI21xp33_ASAP7_75t_L     g340(.A1(new_n904_), .A2(new_n906_1_), .B(new_n908_), .Y(new_n916_1_));
  NOR2xp33_ASAP7_75t_L      g341(.A(new_n916_1_), .B(new_n915_), .Y(new_n917_));
  NOR2xp33_ASAP7_75t_L      g342(.A(new_n914_), .B(new_n917_), .Y(new_n918_));
  NOR4xp25_ASAP7_75t_L      g343(.A(new_n918_), .B(new_n913_), .C(new_n765_), .D(new_n901_1_), .Y(new_n919_));
  A2O1A1Ixp33_ASAP7_75t_L   g344(.A1(n328_o2), .A2(n327_o2), .B(new_n781_1_), .C(new_n917_), .Y(new_n920_));
  NAND2xp33_ASAP7_75t_L     g345(.A(new_n902_), .B(new_n912_), .Y(new_n921_1_));
  NOR2xp33_ASAP7_75t_L      g346(.A(new_n765_), .B(new_n901_1_), .Y(new_n922_));
  AOI21xp33_ASAP7_75t_L     g347(.A1(new_n920_), .A2(new_n921_1_), .B(new_n922_), .Y(new_n923_));
  NOR2xp33_ASAP7_75t_L      g348(.A(new_n923_), .B(new_n919_), .Y(n701));
  AOI21xp33_ASAP7_75t_L     g349(.A1(n276_o2), .A2(n283_o2), .B(n281_o2), .Y(new_n925_));
  INVx1_ASAP7_75t_L         g350(.A(new_n925_), .Y(new_n926_1_));
  NAND2xp33_ASAP7_75t_L     g351(.A(n293_o2), .B(n292_o2), .Y(new_n927_));
  NOR2xp33_ASAP7_75t_L      g352(.A(n293_o2), .B(n292_o2), .Y(new_n928_));
  INVx1_ASAP7_75t_L         g353(.A(new_n928_), .Y(new_n929_));
  NAND3xp33_ASAP7_75t_L     g354(.A(new_n926_1_), .B(new_n929_), .C(new_n927_), .Y(new_n930_));
  INVx1_ASAP7_75t_L         g355(.A(new_n927_), .Y(new_n931_1_));
  OAI21xp33_ASAP7_75t_L     g356(.A1(new_n928_), .A2(new_n931_1_), .B(new_n925_), .Y(new_n932_));
  NAND2xp33_ASAP7_75t_L     g357(.A(new_n932_), .B(new_n930_), .Y(new_n933_));
  NAND2xp33_ASAP7_75t_L     g358(.A(n482_lo_buf_o2), .B(n608_lo_buf_o2), .Y(new_n934_));
  INVx1_ASAP7_75t_L         g359(.A(new_n934_), .Y(new_n935_));
  XNOR2x2_ASAP7_75t_L       g360(.A(new_n935_), .B(new_n933_), .Y(new_n936_1_));
  AND2x2_ASAP7_75t_L        g361(.A(new_n936_1_), .B(n626), .Y(n711));
  NOR2xp33_ASAP7_75t_L      g362(.A(new_n849_), .B(new_n836_1_), .Y(n716));
  AND2x2_ASAP7_75t_L        g363(.A(n1573_o2), .B(n659_lo_buf_o2), .Y(n721));
  NOR3xp33_ASAP7_75t_L      g364(.A(new_n884_), .B(new_n856_1_), .C(new_n885_), .Y(new_n940_));
  AOI21xp33_ASAP7_75t_L     g365(.A1(new_n859_), .A2(new_n882_), .B(new_n858_), .Y(new_n941_1_));
  NAND2xp33_ASAP7_75t_L     g366(.A(n1497_o2), .B(n659_lo_buf_o2), .Y(new_n942_));
  NOR3xp33_ASAP7_75t_L      g367(.A(new_n940_), .B(new_n941_1_), .C(new_n942_), .Y(new_n943_));
  OAI21xp33_ASAP7_75t_L     g368(.A1(new_n941_1_), .A2(new_n940_), .B(new_n942_), .Y(new_n944_));
  A2O1A1O1Ixp25_ASAP7_75t_L g369(.A1(new_n845_), .A2(new_n847_), .B(new_n840_), .C(new_n944_), .D(new_n943_), .Y(n726));
  O2A1O1Ixp33_ASAP7_75t_L   g370(.A1(new_n862_), .A2(new_n864_), .B(new_n869_), .C(new_n897_), .Y(new_n946_1_));
  AOI221xp5_ASAP7_75t_L     g371(.A1(new_n870_), .A2(new_n868_), .B1(new_n892_), .B2(new_n896_1_), .C(new_n863_), .Y(new_n947_));
  NAND2xp33_ASAP7_75t_L     g372(.A(n1625_o2), .B(n647_lo_buf_o2), .Y(new_n948_));
  NOR3xp33_ASAP7_75t_L      g373(.A(new_n946_1_), .B(new_n947_), .C(new_n948_), .Y(new_n949_));
  OAI21xp33_ASAP7_75t_L     g374(.A1(new_n947_), .A2(new_n946_1_), .B(new_n948_), .Y(new_n950_));
  A2O1A1O1Ixp25_ASAP7_75t_L g375(.A1(new_n886_1_), .A2(new_n888_), .B(new_n873_), .C(new_n950_), .D(new_n949_), .Y(n731));
  AND2x2_ASAP7_75t_L        g376(.A(n661), .B(n641), .Y(n736));
  AOI21xp33_ASAP7_75t_L     g377(.A1(new_n914_), .A2(new_n911_1_), .B(new_n915_), .Y(new_n953_));
  AOI21xp33_ASAP7_75t_L     g378(.A1(new_n903_), .A2(n353_o2), .B(n351_o2), .Y(new_n954_));
  XNOR2x2_ASAP7_75t_L       g379(.A(n387_o2), .B(n386_o2), .Y(new_n955_));
  NOR2xp33_ASAP7_75t_L      g380(.A(new_n954_), .B(new_n955_), .Y(new_n956_1_));
  INVx1_ASAP7_75t_L         g381(.A(n351_o2), .Y(new_n957_));
  OAI21xp33_ASAP7_75t_L     g382(.A1(n340_o2), .A2(new_n905_), .B(new_n957_), .Y(new_n958_));
  NAND2xp33_ASAP7_75t_L     g383(.A(n387_o2), .B(n386_o2), .Y(new_n959_));
  OR2x4_ASAP7_75t_L         g384(.A(n387_o2), .B(n386_o2), .Y(new_n960_));
  AOI21xp33_ASAP7_75t_L     g385(.A1(new_n959_), .A2(new_n960_), .B(new_n958_), .Y(new_n961_1_));
  INVx1_ASAP7_75t_L         g386(.A(n1758_o2), .Y(new_n962_));
  INVx1_ASAP7_75t_L         g387(.A(n632_lo_buf_o2), .Y(new_n963_));
  NOR2xp33_ASAP7_75t_L      g388(.A(new_n962_), .B(new_n963_), .Y(new_n964_));
  INVx1_ASAP7_75t_L         g389(.A(new_n964_), .Y(new_n965_));
  NOR3xp33_ASAP7_75t_L      g390(.A(new_n956_1_), .B(new_n961_1_), .C(new_n965_), .Y(new_n966_1_));
  NAND3xp33_ASAP7_75t_L     g391(.A(new_n958_), .B(new_n959_), .C(new_n960_), .Y(new_n967_));
  NAND2xp33_ASAP7_75t_L     g392(.A(new_n954_), .B(new_n955_), .Y(new_n968_));
  AOI21xp33_ASAP7_75t_L     g393(.A1(new_n967_), .A2(new_n968_), .B(new_n964_), .Y(new_n969_));
  NOR3xp33_ASAP7_75t_L      g394(.A(new_n966_1_), .B(new_n953_), .C(new_n969_), .Y(new_n970_));
  OAI21xp33_ASAP7_75t_L     g395(.A1(new_n916_1_), .A2(new_n902_), .B(new_n909_), .Y(new_n971_));
  NAND3xp33_ASAP7_75t_L     g396(.A(new_n967_), .B(new_n968_), .C(new_n964_), .Y(new_n972_));
  OAI21xp33_ASAP7_75t_L     g397(.A1(new_n961_1_), .A2(new_n956_1_), .B(new_n965_), .Y(new_n973_));
  AOI21xp33_ASAP7_75t_L     g398(.A1(new_n972_), .A2(new_n973_), .B(new_n971_), .Y(new_n974_));
  INVx1_ASAP7_75t_L         g399(.A(n1720_o2), .Y(new_n975_));
  NOR2xp33_ASAP7_75t_L      g400(.A(new_n765_), .B(new_n975_), .Y(new_n976_));
  INVx1_ASAP7_75t_L         g401(.A(new_n976_), .Y(new_n977_));
  NOR3xp33_ASAP7_75t_L      g402(.A(new_n970_), .B(new_n974_), .C(new_n977_), .Y(n741));
  XOR2x2_ASAP7_75t_L        g403(.A(n423_o2), .B(n428_o2), .Y(new_n979_));
  NAND2xp33_ASAP7_75t_L     g404(.A(n542_lo_buf_o2), .B(n617_lo_buf_o2), .Y(new_n980_));
  NOR2xp33_ASAP7_75t_L      g405(.A(new_n980_), .B(new_n979_), .Y(new_n981_));
  NOR2xp33_ASAP7_75t_L      g406(.A(n387_o2), .B(n386_o2), .Y(new_n982_));
  A2O1A1Ixp33_ASAP7_75t_L   g407(.A1(new_n904_), .A2(new_n957_), .B(new_n982_), .C(new_n959_), .Y(new_n983_));
  NAND2xp33_ASAP7_75t_L     g408(.A(new_n980_), .B(new_n979_), .Y(new_n984_));
  AOI21xp33_ASAP7_75t_L     g409(.A1(new_n983_), .A2(new_n984_), .B(new_n981_), .Y(new_n985_));
  INVx1_ASAP7_75t_L         g410(.A(n557_lo_buf_o2), .Y(new_n986_));
  INVx1_ASAP7_75t_L         g411(.A(n423_o2), .Y(new_n987_));
  AOI221xp5_ASAP7_75t_L     g412(.A1(n1722_o2), .A2(n572_lo_buf_o2), .B1(n428_o2), .B2(new_n987_), .C(n426_o2), .Y(new_n988_));
  NOR4xp25_ASAP7_75t_L      g413(.A(new_n988_), .B(new_n774_), .C(new_n775_), .D(new_n986_), .Y(new_n989_));
  OA22x2_ASAP7_75t_L        g414(.A1(new_n988_), .A2(new_n774_), .B1(new_n775_), .B2(new_n986_), .Y(new_n990_));
  NOR3xp33_ASAP7_75t_L      g415(.A(new_n985_), .B(new_n990_), .C(new_n989_), .Y(new_n991_));
  NAND2xp33_ASAP7_75t_L     g416(.A(n428_o2), .B(new_n987_), .Y(new_n992_));
  NAND2xp33_ASAP7_75t_L     g417(.A(n423_o2), .B(new_n772_), .Y(new_n993_));
  AND2x2_ASAP7_75t_L        g418(.A(n542_lo_buf_o2), .B(n617_lo_buf_o2), .Y(new_n994_));
  NAND3xp33_ASAP7_75t_L     g419(.A(new_n992_), .B(new_n993_), .C(new_n994_), .Y(new_n995_));
  AND2x2_ASAP7_75t_L        g420(.A(n387_o2), .B(n386_o2), .Y(new_n996_));
  A2O1A1O1Ixp25_ASAP7_75t_L g421(.A1(new_n903_), .A2(n353_o2), .B(n351_o2), .C(new_n960_), .D(new_n996_), .Y(new_n997_));
  AOI21xp33_ASAP7_75t_L     g422(.A1(new_n992_), .A2(new_n993_), .B(new_n994_), .Y(new_n998_));
  OAI21xp33_ASAP7_75t_L     g423(.A1(new_n998_), .A2(new_n997_), .B(new_n995_), .Y(new_n999_));
  NOR2xp33_ASAP7_75t_L      g424(.A(new_n774_), .B(new_n988_), .Y(new_n1000_));
  NOR2xp33_ASAP7_75t_L      g425(.A(new_n775_), .B(new_n986_), .Y(new_n1001_));
  NAND2xp33_ASAP7_75t_L     g426(.A(new_n1001_), .B(new_n1000_), .Y(new_n1002_));
  OAI22xp33_ASAP7_75t_L     g427(.A1(new_n988_), .A2(new_n774_), .B1(new_n775_), .B2(new_n986_), .Y(new_n1003_));
  AOI21xp33_ASAP7_75t_L     g428(.A1(new_n1002_), .A2(new_n1003_), .B(new_n999_), .Y(new_n1004_));
  NAND2xp33_ASAP7_75t_L     g429(.A(n542_lo_buf_o2), .B(n632_lo_buf_o2), .Y(new_n1005_));
  NOR3xp33_ASAP7_75t_L      g430(.A(new_n991_), .B(new_n1004_), .C(new_n1005_), .Y(n746));
  A2O1A1O1Ixp25_ASAP7_75t_L g431(.A1(new_n983_), .A2(new_n984_), .B(new_n981_), .C(new_n1003_), .D(new_n989_), .Y(new_n1007_));
  INVx1_ASAP7_75t_L         g432(.A(new_n773_), .Y(new_n1008_));
  A2O1A1O1Ixp25_ASAP7_75t_L g433(.A1(new_n987_), .A2(n428_o2), .B(n426_o2), .C(new_n1008_), .D(new_n777_), .Y(new_n1009_));
  NOR3xp33_ASAP7_75t_L      g434(.A(new_n1007_), .B(n606), .C(new_n1009_), .Y(n751));
  NAND3xp33_ASAP7_75t_L     g435(.A(new_n846_1_), .B(new_n847_), .C(new_n845_), .Y(new_n1011_));
  OAI21xp33_ASAP7_75t_L     g436(.A1(new_n843_), .A2(new_n840_), .B(new_n825_), .Y(new_n1012_));
  AOI21xp33_ASAP7_75t_L     g437(.A1(new_n1012_), .A2(new_n1011_), .B(new_n851_1_), .Y(new_n1013_));
  NOR2xp33_ASAP7_75t_L      g438(.A(new_n1013_), .B(n681), .Y(n756));
  NAND3xp33_ASAP7_75t_L     g439(.A(new_n888_), .B(new_n886_1_), .C(new_n887_), .Y(new_n1015_));
  OAI21xp33_ASAP7_75t_L     g440(.A1(new_n877_), .A2(new_n873_), .B(new_n860_), .Y(new_n1016_));
  INVx1_ASAP7_75t_L         g441(.A(new_n890_), .Y(new_n1017_));
  AOI21xp33_ASAP7_75t_L     g442(.A1(new_n1015_), .A2(new_n1016_), .B(new_n1017_), .Y(new_n1018_));
  NOR2xp33_ASAP7_75t_L      g443(.A(new_n1018_), .B(n686), .Y(n761));
  A2O1A1Ixp33_ASAP7_75t_L   g444(.A1(new_n874_), .A2(new_n869_), .B(new_n897_), .C(new_n892_), .Y(new_n1020_));
  AOI21xp33_ASAP7_75t_L     g445(.A1(n1682_o2), .A2(n647_lo_buf_o2), .B(new_n1020_), .Y(new_n1021_));
  NOR2xp33_ASAP7_75t_L      g446(.A(n691), .B(new_n1021_), .Y(n766));
  AOI21xp33_ASAP7_75t_L     g447(.A1(new_n845_), .A2(new_n847_), .B(new_n840_), .Y(new_n1023_));
  NAND3xp33_ASAP7_75t_L     g448(.A(new_n858_), .B(new_n859_), .C(new_n882_), .Y(new_n1024_));
  OAI21xp33_ASAP7_75t_L     g449(.A1(new_n885_), .A2(new_n856_1_), .B(new_n884_), .Y(new_n1025_));
  INVx1_ASAP7_75t_L         g450(.A(new_n942_), .Y(new_n1026_));
  AOI21xp33_ASAP7_75t_L     g451(.A1(new_n1024_), .A2(new_n1025_), .B(new_n1026_), .Y(new_n1027_));
  NOR3xp33_ASAP7_75t_L      g452(.A(new_n943_), .B(new_n1027_), .C(new_n1023_), .Y(new_n1028_));
  NAND3xp33_ASAP7_75t_L     g453(.A(new_n1024_), .B(new_n1025_), .C(new_n1026_), .Y(new_n1029_));
  OAI21xp33_ASAP7_75t_L     g454(.A1(new_n825_), .A2(new_n843_), .B(new_n846_1_), .Y(new_n1030_));
  AOI21xp33_ASAP7_75t_L     g455(.A1(new_n944_), .A2(new_n1029_), .B(new_n1030_), .Y(new_n1031_));
  NOR2xp33_ASAP7_75t_L      g456(.A(new_n1031_), .B(new_n1028_), .Y(n771));
  AOI21xp33_ASAP7_75t_L     g457(.A1(new_n888_), .A2(new_n886_1_), .B(new_n873_), .Y(new_n1033_));
  A2O1A1Ixp33_ASAP7_75t_L   g458(.A1(new_n879_), .A2(new_n866_1_), .B(new_n864_), .C(new_n869_), .Y(new_n1034_));
  XOR2x2_ASAP7_75t_L        g459(.A(new_n895_), .B(new_n894_), .Y(new_n1035_));
  NAND2xp33_ASAP7_75t_L     g460(.A(new_n1035_), .B(new_n1034_), .Y(new_n1036_));
  NAND2xp33_ASAP7_75t_L     g461(.A(new_n897_), .B(new_n893_), .Y(new_n1037_));
  INVx1_ASAP7_75t_L         g462(.A(new_n948_), .Y(new_n1038_));
  AOI21xp33_ASAP7_75t_L     g463(.A1(new_n1036_), .A2(new_n1037_), .B(new_n1038_), .Y(new_n1039_));
  NOR3xp33_ASAP7_75t_L      g464(.A(new_n1033_), .B(new_n949_), .C(new_n1039_), .Y(new_n1040_));
  NAND3xp33_ASAP7_75t_L     g465(.A(new_n1036_), .B(new_n1037_), .C(new_n1038_), .Y(new_n1041_));
  OAI21xp33_ASAP7_75t_L     g466(.A1(new_n877_), .A2(new_n860_), .B(new_n887_), .Y(new_n1042_));
  AOI21xp33_ASAP7_75t_L     g467(.A1(new_n950_), .A2(new_n1041_), .B(new_n1042_), .Y(new_n1043_));
  NOR2xp33_ASAP7_75t_L      g468(.A(new_n1043_), .B(new_n1040_), .Y(n776));
  INVx1_ASAP7_75t_L         g469(.A(n696), .Y(new_n1045_));
  NOR3xp33_ASAP7_75t_L      g470(.A(new_n919_), .B(new_n923_), .C(new_n1045_), .Y(n781));
  NOR2xp33_ASAP7_75t_L      g471(.A(new_n765_), .B(new_n962_), .Y(n811));
  NOR2xp33_ASAP7_75t_L      g472(.A(new_n986_), .B(new_n963_), .Y(n816));
  NOR2xp33_ASAP7_75t_L      g473(.A(new_n913_), .B(new_n918_), .Y(new_n1049_));
  MAJIxp5_ASAP7_75t_L       g474(.A(new_n1049_), .B(n696), .C(new_n922_), .Y(n821));
  NOR3xp33_ASAP7_75t_L      g475(.A(new_n997_), .B(new_n981_), .C(new_n998_), .Y(new_n1051_));
  AOI21xp33_ASAP7_75t_L     g476(.A1(new_n984_), .A2(new_n995_), .B(new_n983_), .Y(new_n1052_));
  NAND2xp33_ASAP7_75t_L     g477(.A(n527_lo_buf_o2), .B(n632_lo_buf_o2), .Y(new_n1053_));
  NOR3xp33_ASAP7_75t_L      g478(.A(new_n1051_), .B(new_n1052_), .C(new_n1053_), .Y(new_n1054_));
  OAI21xp33_ASAP7_75t_L     g479(.A1(new_n1052_), .A2(new_n1051_), .B(new_n1053_), .Y(new_n1055_));
  A2O1A1O1Ixp25_ASAP7_75t_L g480(.A1(new_n971_), .A2(new_n973_), .B(new_n966_1_), .C(new_n1055_), .D(new_n1054_), .Y(n826));
  AND4x1_ASAP7_75t_L        g481(.A(n548_lo), .B(n563_lo), .C(n587_lo_buf_o2), .D(n602_lo_buf_o2), .Y(n831));
  NAND4xp25_ASAP7_75t_L     g482(.A(n587_lo_buf_o2), .B(n602_lo_buf_o2), .C(n512_lo_buf_o2), .D(n524_lo_buf_o2), .Y(new_n1058_));
  INVx1_ASAP7_75t_L         g483(.A(new_n1058_), .Y(new_n1059_));
  INVx1_ASAP7_75t_L         g484(.A(n281_o2), .Y(new_n1060_));
  A2O1A1Ixp33_ASAP7_75t_L   g485(.A1(new_n786_1_), .A2(new_n1060_), .B(new_n928_), .C(new_n927_), .Y(new_n1061_));
  AO22x1_ASAP7_75t_L        g486(.A1(n587_lo_buf_o2), .A2(n524_lo_buf_o2), .B1(n602_lo_buf_o2), .B2(n512_lo_buf_o2), .Y(new_n1062_));
  AND4x1_ASAP7_75t_L        g487(.A(n587_lo_buf_o2), .B(n602_lo_buf_o2), .C(n533_lo_buf_o2), .D(n524_lo_buf_o2), .Y(new_n1063_));
  AOI22xp33_ASAP7_75t_L     g488(.A1(n587_lo_buf_o2), .A2(n533_lo_buf_o2), .B1(n602_lo_buf_o2), .B2(n524_lo_buf_o2), .Y(new_n1064_));
  NOR2xp33_ASAP7_75t_L      g489(.A(new_n1064_), .B(new_n1063_), .Y(new_n1065_));
  A2O1A1Ixp33_ASAP7_75t_L   g490(.A1(new_n1061_), .A2(new_n1062_), .B(new_n1059_), .C(new_n1065_), .Y(new_n1066_));
  A2O1A1O1Ixp25_ASAP7_75t_L g491(.A1(new_n929_), .A2(new_n926_1_), .B(new_n931_1_), .C(new_n1062_), .D(new_n1059_), .Y(new_n1067_));
  OAI21xp33_ASAP7_75t_L     g492(.A1(new_n1063_), .A2(new_n1064_), .B(new_n1067_), .Y(new_n1068_));
  AND4x1_ASAP7_75t_L        g493(.A(n512_lo_buf_o2), .B(new_n1068_), .C(n608_lo_buf_o2), .D(new_n1066_), .Y(n836));
  NAND3xp33_ASAP7_75t_L     g494(.A(new_n972_), .B(new_n973_), .C(new_n971_), .Y(new_n1070_));
  OAI21xp33_ASAP7_75t_L     g495(.A1(new_n969_), .A2(new_n966_1_), .B(new_n953_), .Y(new_n1071_));
  AOI21xp33_ASAP7_75t_L     g496(.A1(new_n1071_), .A2(new_n1070_), .B(new_n976_), .Y(new_n1072_));
  NOR2xp33_ASAP7_75t_L      g497(.A(new_n1072_), .B(n741), .Y(n846));
  NAND3xp33_ASAP7_75t_L     g498(.A(new_n1002_), .B(new_n999_), .C(new_n1003_), .Y(new_n1074_));
  OAI21xp33_ASAP7_75t_L     g499(.A1(new_n989_), .A2(new_n990_), .B(new_n985_), .Y(new_n1075_));
  INVx1_ASAP7_75t_L         g500(.A(new_n1005_), .Y(new_n1076_));
  AOI21xp33_ASAP7_75t_L     g501(.A1(new_n1074_), .A2(new_n1075_), .B(new_n1076_), .Y(new_n1077_));
  NOR2xp33_ASAP7_75t_L      g502(.A(new_n1077_), .B(n746), .Y(n851));
  AOI21xp33_ASAP7_75t_L     g503(.A1(new_n971_), .A2(new_n973_), .B(new_n966_1_), .Y(new_n1079_));
  NAND3xp33_ASAP7_75t_L     g504(.A(new_n983_), .B(new_n984_), .C(new_n995_), .Y(new_n1080_));
  OAI21xp33_ASAP7_75t_L     g505(.A1(new_n998_), .A2(new_n981_), .B(new_n997_), .Y(new_n1081_));
  INVx1_ASAP7_75t_L         g506(.A(new_n1053_), .Y(new_n1082_));
  AOI21xp33_ASAP7_75t_L     g507(.A1(new_n1080_), .A2(new_n1081_), .B(new_n1082_), .Y(new_n1083_));
  NOR3xp33_ASAP7_75t_L      g508(.A(new_n1054_), .B(new_n1083_), .C(new_n1079_), .Y(new_n1084_));
  NAND3xp33_ASAP7_75t_L     g509(.A(new_n1080_), .B(new_n1081_), .C(new_n1082_), .Y(new_n1085_));
  OAI21xp33_ASAP7_75t_L     g510(.A1(new_n969_), .A2(new_n953_), .B(new_n972_), .Y(new_n1086_));
  AOI21xp33_ASAP7_75t_L     g511(.A1(new_n1055_), .A2(new_n1085_), .B(new_n1086_), .Y(new_n1087_));
  NOR2xp33_ASAP7_75t_L      g512(.A(new_n1087_), .B(new_n1084_), .Y(n856));
  OA21x2_ASAP7_75t_L        g513(.A1(n606), .A2(new_n1009_), .B(new_n1007_), .Y(new_n1089_));
  NOR2xp33_ASAP7_75t_L      g514(.A(n751), .B(new_n1089_), .Y(n861));
  AND2x2_ASAP7_75t_L        g515(.A(n623_lo), .B(n482_lo_buf_o2), .Y(n871));
  AND2x2_ASAP7_75t_L        g516(.A(n608_lo_buf_o2), .B(n524_lo_buf_o2), .Y(n876));
  NOR2xp33_ASAP7_75t_L      g517(.A(n626), .B(new_n936_1_), .Y(n881));
  NAND3xp33_ASAP7_75t_L     g518(.A(new_n1061_), .B(new_n1058_), .C(new_n1062_), .Y(new_n1094_));
  INVx1_ASAP7_75t_L         g519(.A(new_n1094_), .Y(new_n1095_));
  AOI21xp33_ASAP7_75t_L     g520(.A1(new_n1058_), .A2(new_n1062_), .B(new_n1061_), .Y(new_n1096_));
  NAND2xp33_ASAP7_75t_L     g521(.A(n497_lo_buf_o2), .B(n608_lo_buf_o2), .Y(new_n1097_));
  NOR3xp33_ASAP7_75t_L      g522(.A(new_n1095_), .B(new_n1096_), .C(new_n1097_), .Y(new_n1098_));
  NOR3xp33_ASAP7_75t_L      g523(.A(new_n931_1_), .B(new_n925_), .C(new_n928_), .Y(new_n1099_));
  AOI21xp33_ASAP7_75t_L     g524(.A1(new_n927_), .A2(new_n929_), .B(new_n926_1_), .Y(new_n1100_));
  NOR2xp33_ASAP7_75t_L      g525(.A(new_n1099_), .B(new_n1100_), .Y(new_n1101_));
  MAJIxp5_ASAP7_75t_L       g526(.A(new_n1101_), .B(n626), .C(new_n935_), .Y(new_n1102_));
  AO21x2_ASAP7_75t_L        g527(.A1(new_n1058_), .A2(new_n1062_), .B(new_n1061_), .Y(new_n1103_));
  INVx1_ASAP7_75t_L         g528(.A(new_n1097_), .Y(new_n1104_));
  AOI21xp33_ASAP7_75t_L     g529(.A1(new_n1103_), .A2(new_n1094_), .B(new_n1104_), .Y(new_n1105_));
  NOR3xp33_ASAP7_75t_L      g530(.A(new_n1098_), .B(new_n1102_), .C(new_n1105_), .Y(new_n1106_));
  NOR2xp33_ASAP7_75t_L      g531(.A(new_n1098_), .B(new_n1106_), .Y(n886));
  INVx1_ASAP7_75t_L         g532(.A(new_n1066_), .Y(new_n1108_));
  AND4x1_ASAP7_75t_L        g533(.A(n548_lo), .B(n587_lo_buf_o2), .C(n602_lo_buf_o2), .D(n533_lo_buf_o2), .Y(new_n1109_));
  AOI22xp33_ASAP7_75t_L     g534(.A1(n548_lo), .A2(n587_lo_buf_o2), .B1(n602_lo_buf_o2), .B2(n533_lo_buf_o2), .Y(new_n1110_));
  NOR2xp33_ASAP7_75t_L      g535(.A(new_n1110_), .B(new_n1109_), .Y(new_n1111_));
  O2A1O1Ixp33_ASAP7_75t_L   g536(.A1(new_n1063_), .A2(new_n1108_), .B(new_n1111_), .C(new_n1109_), .Y(n891));
  INVx1_ASAP7_75t_L         g537(.A(a1), .Y(new_n1113_));
  INVx1_ASAP7_75t_L         g538(.A(b0), .Y(new_n1114_));
  NOR2xp33_ASAP7_75t_L      g539(.A(new_n1113_), .B(new_n1114_), .Y(n896));
  INVx1_ASAP7_75t_L         g540(.A(a0), .Y(new_n1116_));
  INVx1_ASAP7_75t_L         g541(.A(b1), .Y(new_n1117_));
  NOR2xp33_ASAP7_75t_L      g542(.A(new_n1116_), .B(new_n1117_), .Y(n901));
  AOI22xp33_ASAP7_75t_L     g543(.A1(n548_lo), .A2(n602_lo_buf_o2), .B1(n563_lo), .B2(n587_lo_buf_o2), .Y(new_n1119_));
  NOR2xp33_ASAP7_75t_L      g544(.A(new_n1119_), .B(n831), .Y(n906));
  AOI22xp33_ASAP7_75t_L     g545(.A1(n512_lo_buf_o2), .A2(n608_lo_buf_o2), .B1(new_n1066_), .B2(new_n1068_), .Y(new_n1121_));
  NOR2xp33_ASAP7_75t_L      g546(.A(new_n1121_), .B(n836), .Y(n911));
  NAND3xp33_ASAP7_75t_L     g547(.A(new_n1103_), .B(new_n1094_), .C(new_n1104_), .Y(new_n1123_));
  INVx1_ASAP7_75t_L         g548(.A(n626), .Y(new_n1124_));
  MAJIxp5_ASAP7_75t_L       g549(.A(new_n933_), .B(new_n934_), .C(new_n1124_), .Y(new_n1125_));
  OAI21xp33_ASAP7_75t_L     g550(.A1(new_n1096_), .A2(new_n1095_), .B(new_n1097_), .Y(new_n1126_));
  AOI21xp33_ASAP7_75t_L     g551(.A1(new_n1126_), .A2(new_n1123_), .B(new_n1125_), .Y(new_n1127_));
  NOR2xp33_ASAP7_75t_L      g552(.A(new_n1106_), .B(new_n1127_), .Y(n916));
  A2O1A1O1Ixp25_ASAP7_75t_L g553(.A1(new_n1062_), .A2(new_n1061_), .B(new_n1059_), .C(new_n1065_), .D(new_n1063_), .Y(new_n1129_));
  XNOR2x2_ASAP7_75t_L       g554(.A(new_n1111_), .B(new_n1129_), .Y(n921));
  INVx1_ASAP7_75t_L         g555(.A(a2), .Y(new_n1131_));
  NOR4xp25_ASAP7_75t_L      g556(.A(new_n1113_), .B(new_n1131_), .C(new_n1114_), .D(new_n1117_), .Y(n931));
  NOR2xp33_ASAP7_75t_L      g557(.A(new_n1131_), .B(new_n1117_), .Y(n946));
  AND2x2_ASAP7_75t_L        g558(.A(a3), .B(b0), .Y(n951));
  NOR4xp25_ASAP7_75t_L      g559(.A(new_n1116_), .B(new_n1113_), .C(new_n1114_), .D(new_n1117_), .Y(n956));
  AOI22xp33_ASAP7_75t_L     g560(.A1(a1), .A2(b1), .B1(a2), .B2(b0), .Y(new_n1136_));
  NOR2xp33_ASAP7_75t_L      g561(.A(new_n1136_), .B(n931), .Y(n966));
  HB1xp67_ASAP7_75t_L       g562(.A(n1221_o2), .Y(n66));
  HB1xp67_ASAP7_75t_L       g563(.A(n1302_o2), .Y(n71));
  HB1xp67_ASAP7_75t_L       g564(.A(a6), .Y(n76));
  HB1xp67_ASAP7_75t_L       g565(.A(n1326_o2), .Y(n81));
  HB1xp67_ASAP7_75t_L       g566(.A(a7), .Y(n86));
  HB1xp67_ASAP7_75t_L       g567(.A(n1368_o2), .Y(n91));
  HB1xp67_ASAP7_75t_L       g568(.A(n1212_o2), .Y(n96));
  HB1xp67_ASAP7_75t_L       g569(.A(b3), .Y(n101));
  HB1xp67_ASAP7_75t_L       g570(.A(b4), .Y(n106));
  HB1xp67_ASAP7_75t_L       g571(.A(n638_lo), .Y(n111));
  HB1xp67_ASAP7_75t_L       g572(.A(b5), .Y(n116));
  HB1xp67_ASAP7_75t_L       g573(.A(n653_lo), .Y(n121));
  HB1xp67_ASAP7_75t_L       g574(.A(b6), .Y(n126));
  HB1xp67_ASAP7_75t_L       g575(.A(n668_lo), .Y(n131));
  HB1xp67_ASAP7_75t_L       g576(.A(n671_lo), .Y(n136));
  HB1xp67_ASAP7_75t_L       g577(.A(b7), .Y(n141));
  HB1xp67_ASAP7_75t_L       g578(.A(n683_lo), .Y(n146));
  HB1xp67_ASAP7_75t_L       g579(.A(n686_lo), .Y(n151));
  HB1xp67_ASAP7_75t_L       g580(.A(n689_lo), .Y(n156));
  HB1xp67_ASAP7_75t_L       g581(.A(n692_lo), .Y(n161));
  HB1xp67_ASAP7_75t_L       g582(.A(n1229_o2), .Y(n166));
  HB1xp67_ASAP7_75t_L       g583(.A(n1228_o2), .Y(n171));
  HB1xp67_ASAP7_75t_L       g584(.A(n1259_o2), .Y(n176));
  HB1xp67_ASAP7_75t_L       g585(.A(n1324_o2), .Y(n181));
  HB1xp67_ASAP7_75t_L       g586(.A(n1325_o2), .Y(n186));
  HB1xp67_ASAP7_75t_L       g587(.A(n1357_o2), .Y(n191));
  HB1xp67_ASAP7_75t_L       g588(.A(n1448_o2), .Y(n196));
  HB1xp67_ASAP7_75t_L       g589(.A(n1449_o2), .Y(n201));
  HB1xp67_ASAP7_75t_L       g590(.A(n1490_o2), .Y(n206));
  HB1xp67_ASAP7_75t_L       g591(.A(n1605_o2), .Y(n211));
  HB1xp67_ASAP7_75t_L       g592(.A(n1609_o2), .Y(n216));
  HB1xp67_ASAP7_75t_L       g593(.A(n1670_o2), .Y(n221));
  HB1xp67_ASAP7_75t_L       g594(.A(n371_o2), .Y(n226));
  HB1xp67_ASAP7_75t_L       g595(.A(n370_o2), .Y(n231));
  HB1xp67_ASAP7_75t_L       g596(.A(n1459_o2), .Y(n236));
  HB1xp67_ASAP7_75t_L       g597(.A(n1460_o2), .Y(n241));
  HB1xp67_ASAP7_75t_L       g598(.A(n1461_o2), .Y(n246));
  HB1xp67_ASAP7_75t_L       g599(.A(n372_o2), .Y(n251));
  HB1xp67_ASAP7_75t_L       g600(.A(n1464_o2), .Y(n256));
  HB1xp67_ASAP7_75t_L       g601(.A(n1497_o2), .Y(n261));
  HB1xp67_ASAP7_75t_L       g602(.A(n1495_o2), .Y(n266));
  HB1xp67_ASAP7_75t_L       g603(.A(n1496_o2), .Y(n271));
  HB1xp67_ASAP7_75t_L       g604(.A(n1520_o2), .Y(n276));
  HB1xp67_ASAP7_75t_L       g605(.A(n1531_o2), .Y(n281));
  HB1xp67_ASAP7_75t_L       g606(.A(n1573_o2), .Y(n286));
  HB1xp67_ASAP7_75t_L       g607(.A(n1625_o2), .Y(n291));
  HB1xp67_ASAP7_75t_L       g608(.A(n1606_o2), .Y(n296));
  HB1xp67_ASAP7_75t_L       g609(.A(n1610_o2), .Y(n301));
  HB1xp67_ASAP7_75t_L       g610(.A(n1635_o2), .Y(n306));
  HB1xp67_ASAP7_75t_L       g611(.A(n415_o2), .Y(n311));
  HB1xp67_ASAP7_75t_L       g612(.A(n1682_o2), .Y(n316));
  HB1xp67_ASAP7_75t_L       g613(.A(n414_o2), .Y(n321));
  HB1xp67_ASAP7_75t_L       g614(.A(n416_o2), .Y(n326));
  HB1xp67_ASAP7_75t_L       g615(.A(n307_o2), .Y(n331));
  HB1xp67_ASAP7_75t_L       g616(.A(n306_o2), .Y(n336));
  HB1xp67_ASAP7_75t_L       g617(.A(n308_o2), .Y(n341));
  HB1xp67_ASAP7_75t_L       g618(.A(n1719_o2), .Y(n346));
  HB1xp67_ASAP7_75t_L       g619(.A(n1720_o2), .Y(n351));
  HB1xp67_ASAP7_75t_L       g620(.A(n1721_o2), .Y(n356));
  HB1xp67_ASAP7_75t_L       g621(.A(n1743_o2), .Y(n361));
  HB1xp67_ASAP7_75t_L       g622(.A(n1751_o2), .Y(n366));
  HB1xp67_ASAP7_75t_L       g623(.A(n1752_o2), .Y(n371));
  HB1xp67_ASAP7_75t_L       g624(.A(n1758_o2), .Y(n376));
  HB1xp67_ASAP7_75t_L       g625(.A(n335_o2), .Y(n381));
  HB1xp67_ASAP7_75t_L       g626(.A(n334_o2), .Y(n386));
  HB1xp67_ASAP7_75t_L       g627(.A(n1765_o2), .Y(n391));
  HB1xp67_ASAP7_75t_L       g628(.A(n527_lo_buf_o2), .Y(n396));
  HB1xp67_ASAP7_75t_L       g629(.A(n336_o2), .Y(n401));
  HB1xp67_ASAP7_75t_L       g630(.A(n542_lo_buf_o2), .Y(n416));
  HB1xp67_ASAP7_75t_L       g631(.A(n287_o2), .Y(n421));
  HB1xp67_ASAP7_75t_L       g632(.A(n286_o2), .Y(n426));
  HB1xp67_ASAP7_75t_L       g633(.A(n557_lo_buf_o2), .Y(n431));
  HB1xp67_ASAP7_75t_L       g634(.A(n659_lo_buf_o2), .Y(n436));
  HB1xp67_ASAP7_75t_L       g635(.A(n288_o2), .Y(n451));
  HB1xp67_ASAP7_75t_L       g636(.A(n572_lo_buf_o2), .Y(n456));
  HB1xp67_ASAP7_75t_L       g637(.A(n632_lo_buf_o2), .Y(n476));
  HB1xp67_ASAP7_75t_L       g638(.A(n482_lo_buf_o2), .Y(n496));
  HB1xp67_ASAP7_75t_L       g639(.A(n497_lo_buf_o2), .Y(n501));
  HB1xp67_ASAP7_75t_L       g640(.A(n587_lo_buf_o2), .Y(n506));
  HB1xp67_ASAP7_75t_L       g641(.A(n602_lo_buf_o2), .Y(n511));
  HB1xp67_ASAP7_75t_L       g642(.A(n467_lo_buf_o2), .Y(n516));
  HB1xp67_ASAP7_75t_L       g643(.A(n274_o2), .Y(n536));
  HB1xp67_ASAP7_75t_L       g644(.A(n275_o2), .Y(n541));
  HB1xp67_ASAP7_75t_L       g645(.A(n512_lo_buf_o2), .Y(n546));
  HB1xp67_ASAP7_75t_L       g646(.A(n276_o2), .Y(n551));
  HB1xp67_ASAP7_75t_L       g647(.A(n524_lo_buf_o2), .Y(n556));
  HB1xp67_ASAP7_75t_L       g648(.A(n674_lo), .Y(n561));
  HB1xp67_ASAP7_75t_L       g649(.A(n641_lo), .Y(n581));
  HB1xp67_ASAP7_75t_L       g650(.A(n533_lo_buf_o2), .Y(n586));
  HB1xp67_ASAP7_75t_L       g651(.A(n608_lo_buf_o2), .Y(n591));
  HB1xp67_ASAP7_75t_L       g652(.A(n548_lo), .Y(n621));
  HB1xp67_ASAP7_75t_L       g653(.A(n563_lo), .Y(n706));
  HB1xp67_ASAP7_75t_L       g654(.A(a1), .Y(n786));
  HB1xp67_ASAP7_75t_L       g655(.A(a2), .Y(n791));
  HB1xp67_ASAP7_75t_L       g656(.A(b0), .Y(n796));
  HB1xp67_ASAP7_75t_L       g657(.A(b1), .Y(n801));
  HB1xp67_ASAP7_75t_L       g658(.A(n656_lo), .Y(n806));
  HB1xp67_ASAP7_75t_L       g659(.A(n623_lo), .Y(n841));
  HB1xp67_ASAP7_75t_L       g660(.A(a0), .Y(n866));
  HB1xp67_ASAP7_75t_L       g661(.A(a3), .Y(n926));
  HB1xp67_ASAP7_75t_L       g662(.A(a5), .Y(n936));
  HB1xp67_ASAP7_75t_L       g663(.A(b2), .Y(n941));
  HB1xp67_ASAP7_75t_L       g664(.A(a4), .Y(n961));
  always @ (posedge clock) begin
    n470_lo <= n66;
    n545_lo <= n71;
    n548_lo <= n76;
    n560_lo <= n81;
    n563_lo <= n86;
    n575_lo <= n91;
    n590_lo <= n96;
    n623_lo <= n101;
    n638_lo <= n106;
    n641_lo <= n111;
    n653_lo <= n116;
    n656_lo <= n121;
    n668_lo <= n126;
    n671_lo <= n131;
    n674_lo <= n136;
    n683_lo <= n141;
    n686_lo <= n146;
    n689_lo <= n151;
    n692_lo <= n156;
    n695_lo <= n161;
    n1001_o2 <= n166;
    n996_o2 <= n171;
    n1011_o2 <= n176;
    n1056_o2 <= n181;
    n1059_o2 <= n186;
    n1074_o2 <= n191;
    n1134_o2 <= n196;
    n1135_o2 <= n201;
    n1158_o2 <= n206;
    n1237_o2 <= n211;
    n1244_o2 <= n216;
    n1266_o2 <= n221;
    n1393_o2 <= n226;
    n1394_o2 <= n231;
    n1210_o2 <= n236;
    n1211_o2 <= n241;
    n1212_o2 <= n246;
    n1437_o2 <= n251;
    n1221_o2 <= n256;
    n1230_o2 <= n261;
    n1228_o2 <= n266;
    n1229_o2 <= n271;
    n1259_o2 <= n276;
    n1265_o2 <= n281;
    n1302_o2 <= n286;
    n1326_o2 <= n291;
    n1324_o2 <= n296;
    n1325_o2 <= n301;
    n1357_o2 <= n306;
    n1648_o2 <= n311;
    n1368_o2 <= n316;
    n1654_o2 <= n321;
    n1700_o2 <= n326;
    n1448_o2 <= n331;
    n1449_o2 <= n336;
    n1490_o2 <= n341;
    n1459_o2 <= n346;
    n1460_o2 <= n351;
    n1461_o2 <= n356;
    n1464_o2 <= n361;
    n1495_o2 <= n366;
    n1496_o2 <= n371;
    n1497_o2 <= n376;
    n1605_o2 <= n381;
    n1609_o2 <= n386;
    n1520_o2 <= n391;
    n1531_o2 <= n396;
    n1670_o2 <= n401;
    n467_o2 <= n406;
    n466_o2 <= n411;
    n1573_o2 <= n416;
    n1606_o2 <= n421;
    n1610_o2 <= n426;
    n1625_o2 <= n431;
    n662_lo_buf_o2 <= n436;
    n468_o2 <= n441;
    n519_o2 <= n446;
    n1635_o2 <= n451;
    n1682_o2 <= n456;
    n371_o2 <= n461;
    n370_o2 <= n466;
    n520_o2 <= n471;
    n1738_o2 <= n476;
    n372_o2 <= n481;
    n307_o2 <= n486;
    n306_o2 <= n491;
    n1719_o2 <= n496;
    n1720_o2 <= n501;
    n1721_o2 <= n506;
    n1722_o2 <= n511;
    n1743_o2 <= n516;
    n523_o2 <= n521;
    n567_o2 <= n526;
    n308_o2 <= n531;
    n1751_o2 <= n536;
    n1752_o2 <= n541;
    n1758_o2 <= n546;
    n1765_o2 <= n551;
    n527_lo_buf_o2 <= n556;
    n677_lo_buf_o2 <= n561;
    n606_o2 <= n566;
    n657_o2 <= n571;
    n568_o2 <= n576;
    n647_lo_buf_o2 <= n581;
    n542_lo_buf_o2 <= n586;
    n617_lo_buf_o2 <= n591;
    n335_o2 <= n596;
    n287_o2 <= n601;
    n530_o2 <= n606;
    n334_o2 <= n611;
    n286_o2 <= n616;
    n557_lo_buf_o2 <= n621;
    n288_o2 <= n626;
    n638_1_o2 <= n631;
    n673_o2 <= n636;
    n415_o2 <= n641;
    n672_o2 <= n646;
    n571_o2 <= n651;
    n646_o2 <= n656;
    n414_o2 <= n661;
    n608_o2 <= n666;
    n659_o2 <= n671;
    n637_o2 <= n676;
    n461_o2 <= n681;
    n551_o2 <= n686;
    n618_o2 <= n691;
    n336_o2 <= n696;
    n367_o2 <= n701;
    n572_lo_buf_o2 <= n706;
    n304_o2 <= n711;
    n509_o2 <= n716;
    n591_o2 <= n721;
    n525_o2 <= n726;
    n615_o2 <= n731;
    n416_o2 <= n736;
    n402_o2 <= n741;
    n489_o2 <= n746;
    n533_o2 <= n751;
    n463_o2 <= n756;
    n553_o2 <= n761;
    n620_o2 <= n766;
    n508_o2 <= n771;
    n590_1_o2 <= n776;
    n368_o2 <= n781;
    n482_lo_buf_o2 <= n786;
    n497_lo_buf_o2 <= n791;
    n587_lo_buf_o2 <= n796;
    n602_lo_buf_o2 <= n801;
    n659_lo_buf_o2 <= n806;
    n446_o2 <= n811;
    n536_o2 <= n816;
    n375_o2 <= n821;
    n474_o2 <= n826;
    n426_o2 <= n831;
    n351_o2 <= n836;
    n632_lo_buf_o2 <= n841;
    n404_o2 <= n846;
    n491_o2 <= n851;
    n445_o2 <= n856;
    n535_o2 <= n861;
    n467_lo_buf_o2 <= n866;
    n328_o2 <= n871;
    n387_o2 <= n876;
    n305_o2 <= n881;
    n340_o2 <= n886;
    n423_o2 <= n891;
    n274_o2 <= n896;
    n275_o2 <= n901;
    n428_o2 <= n906;
    n353_o2 <= n911;
    n327_o2 <= n916;
    n386_o2 <= n921;
    n512_lo_buf_o2 <= n926;
    n281_o2 <= n931;
    n533_lo_buf_o2 <= n936;
    n608_lo_buf_o2 <= n941;
    n293_o2 <= n946;
    n292_o2 <= n951;
    n276_o2 <= n956;
    n524_lo_buf_o2 <= n961;
    n283_o2 <= n966;
  end
  initial begin
    n470_lo <= 1'b0;
    n545_lo <= 1'b0;
    n548_lo <= 1'b0;
    n560_lo <= 1'b0;
    n563_lo <= 1'b0;
    n575_lo <= 1'b0;
    n590_lo <= 1'b0;
    n623_lo <= 1'b0;
    n638_lo <= 1'b0;
    n641_lo <= 1'b0;
    n653_lo <= 1'b0;
    n656_lo <= 1'b0;
    n668_lo <= 1'b0;
    n671_lo <= 1'b0;
    n674_lo <= 1'b0;
    n683_lo <= 1'b0;
    n686_lo <= 1'b0;
    n689_lo <= 1'b0;
    n692_lo <= 1'b0;
    n695_lo <= 1'b0;
    n1001_o2 <= 1'b0;
    n996_o2 <= 1'b0;
    n1011_o2 <= 1'b0;
    n1056_o2 <= 1'b0;
    n1059_o2 <= 1'b0;
    n1074_o2 <= 1'b0;
    n1134_o2 <= 1'b0;
    n1135_o2 <= 1'b0;
    n1158_o2 <= 1'b0;
    n1237_o2 <= 1'b0;
    n1244_o2 <= 1'b0;
    n1266_o2 <= 1'b0;
    n1393_o2 <= 1'b0;
    n1394_o2 <= 1'b0;
    n1210_o2 <= 1'b0;
    n1211_o2 <= 1'b0;
    n1212_o2 <= 1'b0;
    n1437_o2 <= 1'b0;
    n1221_o2 <= 1'b0;
    n1230_o2 <= 1'b0;
    n1228_o2 <= 1'b0;
    n1229_o2 <= 1'b0;
    n1259_o2 <= 1'b0;
    n1265_o2 <= 1'b0;
    n1302_o2 <= 1'b0;
    n1326_o2 <= 1'b0;
    n1324_o2 <= 1'b0;
    n1325_o2 <= 1'b0;
    n1357_o2 <= 1'b0;
    n1648_o2 <= 1'b0;
    n1368_o2 <= 1'b0;
    n1654_o2 <= 1'b0;
    n1700_o2 <= 1'b0;
    n1448_o2 <= 1'b0;
    n1449_o2 <= 1'b0;
    n1490_o2 <= 1'b0;
    n1459_o2 <= 1'b0;
    n1460_o2 <= 1'b0;
    n1461_o2 <= 1'b0;
    n1464_o2 <= 1'b0;
    n1495_o2 <= 1'b0;
    n1496_o2 <= 1'b0;
    n1497_o2 <= 1'b0;
    n1605_o2 <= 1'b0;
    n1609_o2 <= 1'b0;
    n1520_o2 <= 1'b0;
    n1531_o2 <= 1'b0;
    n1670_o2 <= 1'b0;
    n467_o2 <= 1'b0;
    n466_o2 <= 1'b0;
    n1573_o2 <= 1'b0;
    n1606_o2 <= 1'b0;
    n1610_o2 <= 1'b0;
    n1625_o2 <= 1'b0;
    n662_lo_buf_o2 <= 1'b0;
    n468_o2 <= 1'b0;
    n519_o2 <= 1'b0;
    n1635_o2 <= 1'b0;
    n1682_o2 <= 1'b0;
    n371_o2 <= 1'b0;
    n370_o2 <= 1'b0;
    n520_o2 <= 1'b0;
    n1738_o2 <= 1'b0;
    n372_o2 <= 1'b0;
    n307_o2 <= 1'b0;
    n306_o2 <= 1'b0;
    n1719_o2 <= 1'b0;
    n1720_o2 <= 1'b0;
    n1721_o2 <= 1'b0;
    n1722_o2 <= 1'b0;
    n1743_o2 <= 1'b0;
    n523_o2 <= 1'b1;
    n567_o2 <= 1'b0;
    n308_o2 <= 1'b0;
    n1751_o2 <= 1'b0;
    n1752_o2 <= 1'b0;
    n1758_o2 <= 1'b0;
    n1765_o2 <= 1'b0;
    n527_lo_buf_o2 <= 1'b0;
    n677_lo_buf_o2 <= 1'b0;
    n606_o2 <= 1'b0;
    n657_o2 <= 1'b0;
    n568_o2 <= 1'b0;
    n647_lo_buf_o2 <= 1'b0;
    n542_lo_buf_o2 <= 1'b0;
    n617_lo_buf_o2 <= 1'b0;
    n335_o2 <= 1'b0;
    n287_o2 <= 1'b0;
    n530_o2 <= 1'b0;
    n334_o2 <= 1'b0;
    n286_o2 <= 1'b0;
    n557_lo_buf_o2 <= 1'b0;
    n288_o2 <= 1'b0;
    n638_1_o2 <= 1'b0;
    n673_o2 <= 1'b0;
    n415_o2 <= 1'b0;
    n672_o2 <= 1'b1;
    n571_o2 <= 1'b1;
    n646_o2 <= 1'b1;
    n414_o2 <= 1'b0;
    n608_o2 <= 1'b0;
    n659_o2 <= 1'b0;
    n637_o2 <= 1'b0;
    n461_o2 <= 1'b0;
    n551_o2 <= 1'b0;
    n618_o2 <= 1'b0;
    n336_o2 <= 1'b0;
    n367_o2 <= 1'b0;
    n572_lo_buf_o2 <= 1'b0;
    n304_o2 <= 1'b0;
    n509_o2 <= 1'b0;
    n591_o2 <= 1'b0;
    n525_o2 <= 1'b1;
    n615_o2 <= 1'b1;
    n416_o2 <= 1'b0;
    n402_o2 <= 1'b0;
    n489_o2 <= 1'b0;
    n533_o2 <= 1'b0;
    n463_o2 <= 1'b0;
    n553_o2 <= 1'b0;
    n620_o2 <= 1'b0;
    n508_o2 <= 1'b0;
    n590_1_o2 <= 1'b0;
    n368_o2 <= 1'b0;
    n482_lo_buf_o2 <= 1'b0;
    n497_lo_buf_o2 <= 1'b0;
    n587_lo_buf_o2 <= 1'b0;
    n602_lo_buf_o2 <= 1'b0;
    n659_lo_buf_o2 <= 1'b0;
    n446_o2 <= 1'b0;
    n536_o2 <= 1'b0;
    n375_o2 <= 1'b1;
    n474_o2 <= 1'b1;
    n426_o2 <= 1'b0;
    n351_o2 <= 1'b0;
    n632_lo_buf_o2 <= 1'b0;
    n404_o2 <= 1'b0;
    n491_o2 <= 1'b0;
    n445_o2 <= 1'b0;
    n535_o2 <= 1'b0;
    n467_lo_buf_o2 <= 1'b0;
    n328_o2 <= 1'b0;
    n387_o2 <= 1'b0;
    n305_o2 <= 1'b1;
    n340_o2 <= 1'b1;
    n423_o2 <= 1'b1;
    n274_o2 <= 1'b0;
    n275_o2 <= 1'b0;
    n428_o2 <= 1'b0;
    n353_o2 <= 1'b0;
    n327_o2 <= 1'b0;
    n386_o2 <= 1'b0;
    n512_lo_buf_o2 <= 1'b0;
    n281_o2 <= 1'b0;
    n533_lo_buf_o2 <= 1'b0;
    n608_lo_buf_o2 <= 1'b0;
    n293_o2 <= 1'b0;
    n292_o2 <= 1'b0;
    n276_o2 <= 1'b0;
    n524_lo_buf_o2 <= 1'b0;
    n283_o2 <= 1'b0;
  end
endmodule


